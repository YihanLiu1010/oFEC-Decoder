-- HIHO version
-- Take syndrome and hard input data from the syndrome calculator

--library ieee;
--use ieee.std_logic_1164.all;
--
--PACKAGE arr_pkg_9 IS
--    type input_data_array is array (natural range <>) of std_logic_vector(5 downto 0); -- 6 bits
--END; 

library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;
use ieee.math_real.all;
use work.arr_pkg_1.all;
use work.arr_pkg_2.all;
use work.arr_pkg_3.all;

entity bch_decoder_HIHO is
	generic(    
                data_length             : positive := 255;
		input_syndrome_length   : positive := 7;
		softnum     	        : positive := 5 
        );
	port (
		clk             : in std_logic; 					-- system clock
		reset           : in std_logic; 					-- reset
		s1              : in std_logic_vector(7 downto 0);
		s3              : in std_logic_vector(7 downto 0);
		hard_input      : in std_logic_vector(data_length downto 0); 	        -- 6 bits
                soft_input      : in input_data_array(data_length downto 0);
		
		corrections     : out std_logic_vector(2 downto 0);                      -- 100，000，001，010，011
		error_position  : out output_error_location_array(2 downto 0);           -- maximum 3 errors
		hard_output     : out std_logic_vector(data_length downto 0);            -- An array of integer
                soft_output     : out input_data_array(data_length downto 0)
	);
end bch_decoder_HIHO;

architecture rtl of bch_decoder_HIHO is 
-----------------------------------------------------------------------------------------------------------
-- pre-calcaulated array
type table_1 is array (1 to 1275)    of std_logic_vector(7 downto 0);    -- antilog table(255 bits in total)
type table_2 is array (-509 to 1275) of std_logic_vector(1 downto 0);    -- xxxc_1 table
type table_3 is array (0 to 255)     of std_logic_vector(8 downto 0);    -- log table(256 bits in total with one negative number)
type table_4 is array (-509 to 1275) of std_logic_vector(7 downto 0);    -- xxxc_2/3 table
constant log_table      : table_3 := (
        "111111111","000000000","000000001","000011001","000000010","000110010","000011010","011000110","000000011","011011111","000110011","011101110","000011011","001101000","011000111","001001011",
        "000000100","001100100","011100000","000001110","000110100","010001101","011101111","010000001","000011100","011000001","001101001","011111000","011001000","000001000","001001100","001110001",
        "000000101","010001010","001100101","000101111","011100001","000100100","000001111","000100001","000110101","010010011","010001110","011011010","011110000","000010010","010000010","001000101",
        "000011101","010110101","011000010","001111101","001101010","000100111","011111001","010111001","011001001","010011010","000001001","001111000","001001101","011100100","001110010","010100110",
        "000000110","010111111","010001011","001100010","001100110","011011101","000110000","011111101","011100010","010011000","000100101","010110011","000010000","010010001","000100010","010001000",
        "000110110","011010000","010010100","011001110","010001111","010010110","011011011","010111101","011110001","011010010","000010011","001011100","010000011","000111000","001000110","001000000",
        "000011110","001000010","010110110","010100011","011000011","001001000","001111110","001101110","001101011","000111010","000101000","001010100","011111010","010000101","010111010","000111101",
        "011001010","001011110","010011011","010011111","000001010","000010101","001111001","000101011","001001110","011010100","011100101","010101100","001110011","011110011","010100111","001010111",
        "000000111","001110000","011000000","011110111","010001100","010000000","001100011","000001101","001100111","001001010","011011110","011101101","000110001","011000101","011111110","000011000",
        "011100011","010100101","010011001","001110111","000100110","010111000","010110100","001111100","000010001","001000100","010010010","011011001","000100011","000100000","010001001","000101110",
        "000110111","000111111","011010001","001011011","010010101","010111100","011001111","011001101","010010000","010000111","010010111","010110010","011011100","011111100","010111110","001100001",
        "011110010","001010110","011010011","010101011","000010100","000101010","001011101","010011110","010000100","000111100","000111001","001010011","001000111","001101101","001000001","010100010",
        "000011111","000101101","001000011","011011000","010110111","001111011","010100100","001110110","011000100","000010111","001001001","011101100","001111111","000001100","001101111","011110110",
        "001101100","010100001","000111011","001010010","000101001","010011101","001010101","010101010","011111011","001100000","010000110","010110001","010111011","011001100","000111110","001011010",
        "011001011","001011001","001011111","010110000","010011100","010101001","010100000","001010001","000001011","011110101","000010110","011101011","001111010","001110101","000101100","011010111",
        "001001111","010101110","011010101","011101001","011100110","011100111","010101101","011101000","001110100","011010110","011110100","011101010","010101000","001010000","001011000","010101111"
        );
constant antilog_table  : table_1 := (
        "00000001","00000010","00000100","00001000","00010000","00100000","01000000","10000000","00011101","00111010","01110100","11101000","11001101","10000111","00010011","00100110",
        "01001100","10011000","00101101","01011010","10110100","01110101","11101010","11001001","10001111","00000011","00000110","00001100","00011000","00110000","01100000","11000000",
        "10011101","00100111","01001110","10011100","00100101","01001010","10010100","00110101","01101010","11010100","10110101","01110111","11101110","11000001","10011111","00100011",
        "01000110","10001100","00000101","00001010","00010100","00101000","01010000","10100000","01011101","10111010","01101001","11010010","10111001","01101111","11011110","10100001",
        "01011111","10111110","01100001","11000010","10011001","00101111","01011110","10111100","01100101","11001010","10001001","00001111","00011110","00111100","01111000","11110000",
        "11111101","11100111","11010011","10111011","01101011","11010110","10110001","01111111","11111110","11100001","11011111","10100011","01011011","10110110","01110001","11100010",
        "11011001","10101111","01000011","10000110","00010001","00100010","01000100","10001000","00001101","00011010","00110100","01101000","11010000","10111101","01100111","11001110",
        "10000001","00011111","00111110","01111100","11111000","11101101","11000111","10010011","00111011","01110110","11101100","11000101","10010111","00110011","01100110","11001100",
        "10000101","00010111","00101110","01011100","10111000","01101101","11011010","10101001","01001111","10011110","00100001","01000010","10000100","00010101","00101010","01010100",
        "10101000","01001101","10011010","00101001","01010010","10100100","01010101","10101010","01001001","10010010","00111001","01110010","11100100","11010101","10110111","01110011",
        "11100110","11010001","10111111","01100011","11000110","10010001","00111111","01111110","11111100","11100101","11010111","10110011","01111011","11110110","11110001","11111111",
        "11100011","11011011","10101011","01001011","10010110","00110001","01100010","11000100","10010101","00110111","01101110","11011100","10100101","01010111","10101110","01000001",
        "10000010","00011001","00110010","01100100","11001000","10001101","00000111","00001110","00011100","00111000","01110000","11100000","11011101","10100111","01010011","10100110",
        "01010001","10100010","01011001","10110010","01111001","11110010","11111001","11101111","11000011","10011011","00101011","01010110","10101100","01000101","10001010","00001001",
        "00010010","00100100","01001000","10010000","00111101","01111010","11110100","11110101","11110111","11110011","11111011","11101011","11001011","10001011","00001011","00010110",
        "00101100","01011000","10110000","01111101","11111010","11101001","11001111","10000011","00011011","00110110","01101100","11011000","10101101","01000111","10001110",
        "00000001","00000010","00000100","00001000","00010000","00100000","01000000","10000000","00011101","00111010","01110100","11101000","11001101","10000111","00010011","00100110",
        "01001100","10011000","00101101","01011010","10110100","01110101","11101010","11001001","10001111","00000011","00000110","00001100","00011000","00110000","01100000","11000000",
        "10011101","00100111","01001110","10011100","00100101","01001010","10010100","00110101","01101010","11010100","10110101","01110111","11101110","11000001","10011111","00100011",
        "01000110","10001100","00000101","00001010","00010100","00101000","01010000","10100000","01011101","10111010","01101001","11010010","10111001","01101111","11011110","10100001",
        "01011111","10111110","01100001","11000010","10011001","00101111","01011110","10111100","01100101","11001010","10001001","00001111","00011110","00111100","01111000","11110000",
        "11111101","11100111","11010011","10111011","01101011","11010110","10110001","01111111","11111110","11100001","11011111","10100011","01011011","10110110","01110001","11100010",
        "11011001","10101111","01000011","10000110","00010001","00100010","01000100","10001000","00001101","00011010","00110100","01101000","11010000","10111101","01100111","11001110",
        "10000001","00011111","00111110","01111100","11111000","11101101","11000111","10010011","00111011","01110110","11101100","11000101","10010111","00110011","01100110","11001100",
        "10000101","00010111","00101110","01011100","10111000","01101101","11011010","10101001","01001111","10011110","00100001","01000010","10000100","00010101","00101010","01010100",
        "10101000","01001101","10011010","00101001","01010010","10100100","01010101","10101010","01001001","10010010","00111001","01110010","11100100","11010101","10110111","01110011",
        "11100110","11010001","10111111","01100011","11000110","10010001","00111111","01111110","11111100","11100101","11010111","10110011","01111011","11110110","11110001","11111111",
        "11100011","11011011","10101011","01001011","10010110","00110001","01100010","11000100","10010101","00110111","01101110","11011100","10100101","01010111","10101110","01000001",
        "10000010","00011001","00110010","01100100","11001000","10001101","00000111","00001110","00011100","00111000","01110000","11100000","11011101","10100111","01010011","10100110",
        "01010001","10100010","01011001","10110010","01111001","11110010","11111001","11101111","11000011","10011011","00101011","01010110","10101100","01000101","10001010","00001001",
        "00010010","00100100","01001000","10010000","00111101","01111010","11110100","11110101","11110111","11110011","11111011","11101011","11001011","10001011","00001011","00010110",
        "00101100","01011000","10110000","01111101","11111010","11101001","11001111","10000011","00011011","00110110","01101100","11011000","10101101","01000111","10001110",
        "00000001","00000010","00000100","00001000","00010000","00100000","01000000","10000000","00011101","00111010","01110100","11101000","11001101","10000111","00010011","00100110",
        "01001100","10011000","00101101","01011010","10110100","01110101","11101010","11001001","10001111","00000011","00000110","00001100","00011000","00110000","01100000","11000000",
        "10011101","00100111","01001110","10011100","00100101","01001010","10010100","00110101","01101010","11010100","10110101","01110111","11101110","11000001","10011111","00100011",
        "01000110","10001100","00000101","00001010","00010100","00101000","01010000","10100000","01011101","10111010","01101001","11010010","10111001","01101111","11011110","10100001",
        "01011111","10111110","01100001","11000010","10011001","00101111","01011110","10111100","01100101","11001010","10001001","00001111","00011110","00111100","01111000","11110000",
        "11111101","11100111","11010011","10111011","01101011","11010110","10110001","01111111","11111110","11100001","11011111","10100011","01011011","10110110","01110001","11100010",
        "11011001","10101111","01000011","10000110","00010001","00100010","01000100","10001000","00001101","00011010","00110100","01101000","11010000","10111101","01100111","11001110",
        "10000001","00011111","00111110","01111100","11111000","11101101","11000111","10010011","00111011","01110110","11101100","11000101","10010111","00110011","01100110","11001100",
        "10000101","00010111","00101110","01011100","10111000","01101101","11011010","10101001","01001111","10011110","00100001","01000010","10000100","00010101","00101010","01010100",
        "10101000","01001101","10011010","00101001","01010010","10100100","01010101","10101010","01001001","10010010","00111001","01110010","11100100","11010101","10110111","01110011",
        "11100110","11010001","10111111","01100011","11000110","10010001","00111111","01111110","11111100","11100101","11010111","10110011","01111011","11110110","11110001","11111111",
        "11100011","11011011","10101011","01001011","10010110","00110001","01100010","11000100","10010101","00110111","01101110","11011100","10100101","01010111","10101110","01000001",
        "10000010","00011001","00110010","01100100","11001000","10001101","00000111","00001110","00011100","00111000","01110000","11100000","11011101","10100111","01010011","10100110",
        "01010001","10100010","01011001","10110010","01111001","11110010","11111001","11101111","11000011","10011011","00101011","01010110","10101100","01000101","10001010","00001001",
        "00010010","00100100","01001000","10010000","00111101","01111010","11110100","11110101","11110111","11110011","11111011","11101011","11001011","10001011","00001011","00010110",
        "00101100","01011000","10110000","01111101","11111010","11101001","11001111","10000011","00011011","00110110","01101100","11011000","10101101","01000111","10001110",
        "00000001","00000010","00000100","00001000","00010000","00100000","01000000","10000000","00011101","00111010","01110100","11101000","11001101","10000111","00010011","00100110",
        "01001100","10011000","00101101","01011010","10110100","01110101","11101010","11001001","10001111","00000011","00000110","00001100","00011000","00110000","01100000","11000000",
        "10011101","00100111","01001110","10011100","00100101","01001010","10010100","00110101","01101010","11010100","10110101","01110111","11101110","11000001","10011111","00100011",
        "01000110","10001100","00000101","00001010","00010100","00101000","01010000","10100000","01011101","10111010","01101001","11010010","10111001","01101111","11011110","10100001",
        "01011111","10111110","01100001","11000010","10011001","00101111","01011110","10111100","01100101","11001010","10001001","00001111","00011110","00111100","01111000","11110000",
        "11111101","11100111","11010011","10111011","01101011","11010110","10110001","01111111","11111110","11100001","11011111","10100011","01011011","10110110","01110001","11100010",
        "11011001","10101111","01000011","10000110","00010001","00100010","01000100","10001000","00001101","00011010","00110100","01101000","11010000","10111101","01100111","11001110",
        "10000001","00011111","00111110","01111100","11111000","11101101","11000111","10010011","00111011","01110110","11101100","11000101","10010111","00110011","01100110","11001100",
        "10000101","00010111","00101110","01011100","10111000","01101101","11011010","10101001","01001111","10011110","00100001","01000010","10000100","00010101","00101010","01010100",
        "10101000","01001101","10011010","00101001","01010010","10100100","01010101","10101010","01001001","10010010","00111001","01110010","11100100","11010101","10110111","01110011",
        "11100110","11010001","10111111","01100011","11000110","10010001","00111111","01111110","11111100","11100101","11010111","10110011","01111011","11110110","11110001","11111111",
        "11100011","11011011","10101011","01001011","10010110","00110001","01100010","11000100","10010101","00110111","01101110","11011100","10100101","01010111","10101110","01000001",
        "10000010","00011001","00110010","01100100","11001000","10001101","00000111","00001110","00011100","00111000","01110000","11100000","11011101","10100111","01010011","10100110",
        "01010001","10100010","01011001","10110010","01111001","11110010","11111001","11101111","11000011","10011011","00101011","01010110","10101100","01000101","10001010","00001001",
        "00010010","00100100","01001000","10010000","00111101","01111010","11110100","11110101","11110111","11110011","11111011","11101011","11001011","10001011","00001011","00010110",
        "00101100","01011000","10110000","01111101","11111010","11101001","11001111","10000011","00011011","00110110","01101100","11011000","10101101","01000111","10001110",
        "00000001","00000010","00000100","00001000","00010000","00100000","01000000","10000000","00011101","00111010","01110100","11101000","11001101","10000111","00010011","00100110",
        "01001100","10011000","00101101","01011010","10110100","01110101","11101010","11001001","10001111","00000011","00000110","00001100","00011000","00110000","01100000","11000000",
        "10011101","00100111","01001110","10011100","00100101","01001010","10010100","00110101","01101010","11010100","10110101","01110111","11101110","11000001","10011111","00100011",
        "01000110","10001100","00000101","00001010","00010100","00101000","01010000","10100000","01011101","10111010","01101001","11010010","10111001","01101111","11011110","10100001",
        "01011111","10111110","01100001","11000010","10011001","00101111","01011110","10111100","01100101","11001010","10001001","00001111","00011110","00111100","01111000","11110000",
        "11111101","11100111","11010011","10111011","01101011","11010110","10110001","01111111","11111110","11100001","11011111","10100011","01011011","10110110","01110001","11100010",
        "11011001","10101111","01000011","10000110","00010001","00100010","01000100","10001000","00001101","00011010","00110100","01101000","11010000","10111101","01100111","11001110",
        "10000001","00011111","00111110","01111100","11111000","11101101","11000111","10010011","00111011","01110110","11101100","11000101","10010111","00110011","01100110","11001100",
        "10000101","00010111","00101110","01011100","10111000","01101101","11011010","10101001","01001111","10011110","00100001","01000010","10000100","00010101","00101010","01010100",
        "10101000","01001101","10011010","00101001","01010010","10100100","01010101","10101010","01001001","10010010","00111001","01110010","11100100","11010101","10110111","01110011",
        "11100110","11010001","10111111","01100011","11000110","10010001","00111111","01111110","11111100","11100101","11010111","10110011","01111011","11110110","11110001","11111111",
        "11100011","11011011","10101011","01001011","10010110","00110001","01100010","11000100","10010101","00110111","01101110","11011100","10100101","01010111","10101110","01000001",
        "10000010","00011001","00110010","01100100","11001000","10001101","00000111","00001110","00011100","00111000","01110000","11100000","11011101","10100111","01010011","10100110",
        "01010001","10100010","01011001","10110010","01111001","11110010","11111001","11101111","11000011","10011011","00101011","01010110","10101100","01000101","10001010","00001001",
        "00010010","00100100","01001000","10010000","00111101","01111010","11110100","11110101","11110111","11110011","11111011","11101011","11001011","10001011","00001011","00010110",
        "00101100","01011000","10110000","01111101","11111010","11101001","11001111","10000011","00011011","00110110","01101100","11011000","10101101","01000111","10001110");
constant xxxc_1  		: table_2 := (
        "10","10","10","10","10","00","10","10","10","00","00","00","10","10","10","00",
        "10","10","00","10","00","00","00","10","10","10","10","10","10","00","00","10",
        "10","00","10","10","00","10","10","00","00","10","00","00","00","10","10","00",
        "10","10","10","10","10","00","10","00","10","00","00","10","00","00","10","00",
        "10","00","00","10","10","00","10","00","00","10","10","10","10","00","00","00",
        "00","00","10","00","00","10","00","00","00","00","10","00","10","00","00","00",
        "10","00","10","10","10","00","10","10","10","10","00","00","10","00","00","10",
        "10","10","00","00","00","00","10","10","00","00","00","10","10","00","00","10",
        "10","10","00","10","00","00","10","00","10","10","00","10","10","10","00","10",
        "00","10","10","00","10","00","10","00","10","10","00","00","00","10","00","00",
        "00","10","00","00","10","10","00","00","00","00","10","00","00","00","00","00",
        "00","10","00","10","10","00","00","10","10","00","00","10","00","10","00","10",
        "10","10","00","00","10","10","10","10","10","00","00","00","10","00","10","00",
        "10","00","10","00","00","00","00","00","10","10","00","10","00","10","10","10",
        "10","00","10","10","00","00","00","00","00","00","00","00","10","10","10","10",
        "00","10","00","00","00","00","10","10","10","00","00","10","00","10","10",
        "10","10","10","10","10","00","10","10","10","00","00","00","10","10","10","00",
        "10","10","00","10","00","00","00","10","10","10","10","10","10","00","00","10",
        "10","00","10","10","00","10","10","00","00","10","00","00","00","10","10","00",
        "10","10","10","10","10","00","10","00","10","00","00","10","00","00","10","00",
        "10","00","00","10","10","00","10","00","00","10","10","10","10","00","00","00",
        "00","00","10","00","00","10","00","00","00","00","10","00","10","00","00","00",
        "10","00","10","10","10","00","10","10","10","10","00","00","10","00","00","10",
        "10","10","00","00","00","00","10","10","00","00","00","10","10","00","00","10",
        "10","10","00","10","00","00","10","00","10","10","00","10","10","10","00","10",
        "00","10","10","00","10","00","10","00","10","10","00","00","00","10","00","00",
        "00","10","00","00","10","10","00","00","00","00","10","00","00","00","00","00",
        "00","10","00","10","10","00","00","10","10","00","00","10","00","10","00","10",
        "10","10","00","00","10","10","10","10","10","00","00","00","10","00","10","00",
        "10","00","10","00","00","00","00","00","10","10","00","10","00","10","10","10",
        "10","00","10","10","00","00","00","00","00","00","00","00","10","10","10","10",
        "00","10","00","00","00","00","10","10","10","00","00","10","00","10","10",
        "10","10","10","10","10","00","10","10","10","00","00","00","10","10","10","00",
        "10","10","00","10","00","00","00","10","10","10","10","10","10","00","00","10",
        "10","00","10","10","00","10","10","00","00","10","00","00","00","10","10","00",
        "10","10","10","10","10","00","10","00","10","00","00","10","00","00","10","00",
        "10","00","00","10","10","00","10","00","00","10","10","10","10","00","00","00",
        "00","00","10","00","00","10","00","00","00","00","10","00","10","00","00","00",
        "10","00","10","10","10","00","10","10","10","10","00","00","10","00","00","10",
        "10","10","00","00","00","00","10","10","00","00","00","10","10","00","00","10",
        "10","10","00","10","00","00","10","00","10","10","00","10","10","10","00","10",
        "00","10","10","00","10","00","10","00","10","10","00","00","00","10","00","00",
        "00","10","00","00","10","10","00","00","00","00","10","00","00","00","00","00",
        "00","10","00","10","10","00","00","10","10","00","00","10","00","10","00","10",
        "10","10","00","00","10","10","10","10","10","00","00","00","10","00","10","00",
        "10","00","10","00","00","00","00","00","10","10","00","10","00","10","10","10",
        "10","00","10","10","00","00","00","00","00","00","00","00","10","10","10","10",
        "00","10","00","00","00","00","10","10","10","00","00","10","00","10","10",
        "10","10","10","10","10","00","10","10","10","00","00","00","10","10","10","00",
        "10","10","00","10","00","00","00","10","10","10","10","10","10","00","00","10",
        "10","00","10","10","00","10","10","00","00","10","00","00","00","10","10","00",
        "10","10","10","10","10","00","10","00","10","00","00","10","00","00","10","00",
        "10","00","00","10","10","00","10","00","00","10","10","10","10","00","00","00",
        "00","00","10","00","00","10","00","00","00","00","10","00","10","00","00","00",
        "10","00","10","10","10","00","10","10","10","10","00","00","10","00","00","10",
        "10","10","00","00","00","00","10","10","00","00","00","10","10","00","00","10",
        "10","10","00","10","00","00","10","00","10","10","00","10","10","10","00","10",
        "00","10","10","00","10","00","10","00","10","10","00","00","00","10","00","00",
        "00","10","00","00","10","10","00","00","00","00","10","00","00","00","00","00",
        "00","10","00","10","10","00","00","10","10","00","00","10","00","10","00","10",
        "10","10","00","00","10","10","10","10","10","00","00","00","10","00","10","00",
        "10","00","10","00","00","00","00","00","10","10","00","10","00","10","10","10",
        "10","00","10","10","00","00","00","00","00","00","00","00","10","10","10","10",
        "00","10","00","00","00","00","10","10","10","00","00","10","00","10","10",
        "10","10","10","10","10","00","10","10","10","00","00","00","10","10","10","00",
        "10","10","00","10","00","00","00","10","10","10","10","10","10","00","00","10",
        "10","00","10","10","00","10","10","00","00","10","00","00","00","10","10","00",
        "10","10","10","10","10","00","10","00","10","00","00","10","00","00","10","00",
        "10","00","00","10","10","00","10","00","00","10","10","10","10","00","00","00",
        "00","00","10","00","00","10","00","00","00","00","10","00","10","00","00","00",
        "10","00","10","10","10","00","10","10","10","10","00","00","10","00","00","10",
        "10","10","00","00","00","00","10","10","00","00","00","10","10","00","00","10",
        "10","10","00","10","00","00","10","00","10","10","00","10","10","10","00","10",
        "00","10","10","00","10","00","10","00","10","10","00","00","00","10","00","00",
        "00","10","00","00","10","10","00","00","00","00","10","00","00","00","00","00",
        "00","10","00","10","10","00","00","10","10","00","00","10","00","10","00","10",
        "10","10","00","00","10","10","10","10","10","00","00","00","10","00","10","00",
        "10","00","10","00","00","00","00","00","10","10","00","10","00","10","10","10",
        "10","00","10","10","00","00","00","00","00","00","00","00","10","10","10","10",
        "00","10","00","00","00","00","10","10","10","00","00","10","00","10","10",
        "10","10","10","10","10","00","10","10","10","00","00","00","10","10","10","00",
        "10","10","00","10","00","00","00","10","10","10","10","10","10","00","00","10",
        "10","00","10","10","00","10","10","00","00","10","00","00","00","10","10","00",
        "10","10","10","10","10","00","10","00","10","00","00","10","00","00","10","00",
        "10","00","00","10","10","00","10","00","00","10","10","10","10","00","00","00",
        "00","00","10","00","00","10","00","00","00","00","10","00","10","00","00","00",
        "10","00","10","10","10","00","10","10","10","10","00","00","10","00","00","10",
        "10","10","00","00","00","00","10","10","00","00","00","10","10","00","00","10",
        "10","10","00","10","00","00","10","00","10","10","00","10","10","10","00","10",
        "00","10","10","00","10","00","10","00","10","10","00","00","00","10","00","00",
        "00","10","00","00","10","10","00","00","00","00","10","00","00","00","00","00",
        "00","10","00","10","10","00","00","10","10","00","00","10","00","10","00","10",
        "10","10","00","00","10","10","10","10","10","00","00","00","10","00","10","00",
        "10","00","10","00","00","00","00","00","10","10","00","10","00","10","10","10",
        "10","00","10","10","00","00","00","00","00","00","00","00","10","10","10","10",
        "00","10","00","00","00","00","10","10","10","00","00","10","00","10","10",
        "10","10","10","10","10","00","10","10","10","00","00","00","10","10","10","00",
        "10","10","00","10","00","00","00","10","10","10","10","10","10","00","00","10",
        "10","00","10","10","00","10","10","00","00","10","00","00","00","10","10","00",
        "10","10","10","10","10","00","10","00","10","00","00","10","00","00","10","00",
        "10","00","00","10","10","00","10","00","00","10","10","10","10","00","00","00",
        "00","00","10","00","00","10","00","00","00","00","10","00","10","00","00","00",
        "10","00","10","10","10","00","10","10","10","10","00","00","10","00","00","10",
        "10","10","00","00","00","00","10","10","00","00","00","10","10","00","00","10",
        "10","10","00","10","00","00","10","00","10","10","00","10","10","10","00","10",
        "00","10","10","00","10","00","10","00","10","10","00","00","00","10","00","00",
        "00","10","00","00","10","10","00","00","00","00","10","00","00","00","00","00",
        "00","10","00","10","10","00","00","10","10","00","00","10","00","10","00","10",
        "10","10","00","00","10","10","10","10","10","00","00","00","10","00","10","00",
        "10","00","10","00","00","00","00","00","10","10","00","10","00","10","10","10",
        "10","00","10","10","00","00","00","00","00","00","00","00","10","10","10","10",
        "00","10","00","00","00","00","10","10","10","00","00","10","00","10","10");
constant xxxc_2         : table_4 := (
        "01010101","00001011","00010110","00010010","00101100","00000000","00100100","00110110","01011000","00000000","00000000","00000000","01001000","10000000","01101100","00000000",
        "01011111","01110111","00000000","01001011","00000000","00000000","00000000","00011000","10000111","01110010","00000001","01110110","01000011","00000000","00000000","00001010",
        "01100001","00000000","00110011","01001110","00000000","01011001","10001111","00000000","00000000","01011110","00000000","00000000","00000000","01011011","00110000","00000000",
        "00001111","01111100","01001101","01111011","00000010","00000000","01001001","00000000","10000110","00000000","00000000","10011011","00000000","00000000","00010100","00000000",
        "01111101","00000000","00000000","00100000","01100110","00000000","10011100","00000000","00000000","01010110","10010111","01110100","00011111","00000000","00000000","00000000",
        "00000000","00000000","10010101","00000000","00000000","00010001","00000000","00000000","00000000","00000000","10100011","00000000","01100000","00000000","00000000","00000000",
        "00011110","00000000","01101001","10010100","10011010","00000000","01101111","01110011","00000100","10001110","00000000","00000000","10010010","00000000","00000000","00010011",
        "00001101","10000001","00000000","00000000","00000000","00000000","00110111","00000111","00000000","00000000","00000000","10011000","00101000","00000000","00000000","10101011",
        "10000101","00001001","00000000","00011011","00000000","00000000","01000000","00000000","10111011","10100101","00000000","00001100","00111001","00111011","00000000","00000101",
        "00000000","00100111","10101100","00000000","00101111","00000000","10101101","00000000","00111110","10111101","00000000","00000000","00000000","11001101","00000000","00000000",
        "00000000","00010000","00000000","00000000","00101011","00111010","00000000","00000000","00000000","00000000","00100010","00000000","00000000","00000000","00000000","00000000",
        "00000000","01001010","00000000","10111001","01000111","00000000","00000000","00101110","11000000","00000000","00000000","00111000","00000000","01001100","00000000","11010101",
        "00111100","00110100","00000000","00000000","11010010","00000110","00101001","01000101","00110101","00000000","00000000","00000000","11011110","00000000","11100110","00000000",
        "00001000","00000000","00011101","00000000","00000000","00000000","00000000","00000000","00100101","11011100","00000000","00010111","00000000","00011100","00100110","11101010",
        "00011010","00000000","00000011","01000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01101110","01100010","00001110","01110101",
        "00000000","01010001","00000000","00000000","00000000","00000000","00110001","00111101","01010000","00000000","00000000","01011101","00000000","01001111","01010111","01010101",
        "00001011","00010110","00010010","00101100","00000000","00100100","00110110","01011000","00000000","00000000","00000000","01001000","10000000","01101100","00000000","01011111",
        "01110111","00000000","01001011","00000000","00000000","00000000","00011000","10000111","01110010","00000001","01110110","01000011","00000000","00000000","00001010","01100001",
        "00000000","00110011","01001110","00000000","01011001","10001111","00000000","00000000","01011110","00000000","00000000","00000000","01011011","00110000","00000000","00001111",
        "01111100","01001101","01111011","00000010","00000000","01001001","00000000","10000110","00000000","00000000","10011011","00000000","00000000","00010100","00000000","01111101",
        "00000000","00000000","00100000","01100110","00000000","10011100","00000000","00000000","01010110","10010111","01110100","00011111","00000000","00000000","00000000","00000000",
        "00000000","10010101","00000000","00000000","00010001","00000000","00000000","00000000","00000000","10100011","00000000","01100000","00000000","00000000","00000000","00011110",
        "00000000","01101001","10010100","10011010","00000000","01101111","01110011","00000100","10001110","00000000","00000000","10010010","00000000","00000000","00010011","00001101",
        "10000001","00000000","00000000","00000000","00000000","00110111","00000111","00000000","00000000","00000000","10011000","00101000","00000000","00000000","10101011","10000101",
        "00001001","00000000","00011011","00000000","00000000","01000000","00000000","10111011","10100101","00000000","00001100","00111001","00111011","00000000","00000101","00000000",
        "00100111","10101100","00000000","00101111","00000000","10101101","00000000","00111110","10111101","00000000","00000000","00000000","11001101","00000000","00000000","00000000",
        "00010000","00000000","00000000","00101011","00111010","00000000","00000000","00000000","00000000","00100010","00000000","00000000","00000000","00000000","00000000","00000000",
        "01001010","00000000","10111001","01000111","00000000","00000000","00101110","11000000","00000000","00000000","00111000","00000000","01001100","00000000","11010101","00111100",
        "00110100","00000000","00000000","11010010","00000110","00101001","01000101","00110101","00000000","00000000","00000000","11011110","00000000","11100110","00000000","00001000",
        "00000000","00011101","00000000","00000000","00000000","00000000","00000000","00100101","11011100","00000000","00010111","00000000","00011100","00100110","11101010","00011010",
        "00000000","00000011","01000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01101110","01100010","00001110","01110101","00000000",
        "01010001","00000000","00000000","00000000","00000000","00110001","00111101","01010000","00000000","00000000","01011101","00000000","01001111","01010111",
        "01010101","00001011","00010110","00010010","00101100","00000000","00100100","00110110","01011000","00000000","00000000","00000000","01001000","10000000","01101100","00000000",
        "01011111","01110111","00000000","01001011","00000000","00000000","00000000","00011000","10000111","01110010","00000001","01110110","01000011","00000000","00000000","00001010",
        "01100001","00000000","00110011","01001110","00000000","01011001","10001111","00000000","00000000","01011110","00000000","00000000","00000000","01011011","00110000","00000000",
        "00001111","01111100","01001101","01111011","00000010","00000000","01001001","00000000","10000110","00000000","00000000","10011011","00000000","00000000","00010100","00000000",
        "01111101","00000000","00000000","00100000","01100110","00000000","10011100","00000000","00000000","01010110","10010111","01110100","00011111","00000000","00000000","00000000",
        "00000000","00000000","10010101","00000000","00000000","00010001","00000000","00000000","00000000","00000000","10100011","00000000","01100000","00000000","00000000","00000000",
        "00011110","00000000","01101001","10010100","10011010","00000000","01101111","01110011","00000100","10001110","00000000","00000000","10010010","00000000","00000000","00010011",
        "00001101","10000001","00000000","00000000","00000000","00000000","00110111","00000111","00000000","00000000","00000000","10011000","00101000","00000000","00000000","10101011",
        "10000101","00001001","00000000","00011011","00000000","00000000","01000000","00000000","10111011","10100101","00000000","00001100","00111001","00111011","00000000","00000101",
        "00000000","00100111","10101100","00000000","00101111","00000000","10101101","00000000","00111110","10111101","00000000","00000000","00000000","11001101","00000000","00000000",
        "00000000","00010000","00000000","00000000","00101011","00111010","00000000","00000000","00000000","00000000","00100010","00000000","00000000","00000000","00000000","00000000",
        "00000000","01001010","00000000","10111001","01000111","00000000","00000000","00101110","11000000","00000000","00000000","00111000","00000000","01001100","00000000","11010101",
        "00111100","00110100","00000000","00000000","11010010","00000110","00101001","01000101","00110101","00000000","00000000","00000000","11011110","00000000","11100110","00000000",
        "00001000","00000000","00011101","00000000","00000000","00000000","00000000","00000000","00100101","11011100","00000000","00010111","00000000","00011100","00100110","11101010",
        "00011010","00000000","00000011","01000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01101110","01100010","00001110","01110101",
        "00000000","01010001","00000000","00000000","00000000","00000000","00110001","00111101","01010000","00000000","00000000","01011101","00000000","01001111","01010111","01010101",
        "00001011","00010110","00010010","00101100","00000000","00100100","00110110","01011000","00000000","00000000","00000000","01001000","10000000","01101100","00000000","01011111",
        "01110111","00000000","01001011","00000000","00000000","00000000","00011000","10000111","01110010","00000001","01110110","01000011","00000000","00000000","00001010","01100001",
        "00000000","00110011","01001110","00000000","01011001","10001111","00000000","00000000","01011110","00000000","00000000","00000000","01011011","00110000","00000000","00001111",
        "01111100","01001101","01111011","00000010","00000000","01001001","00000000","10000110","00000000","00000000","10011011","00000000","00000000","00010100","00000000","01111101",
        "00000000","00000000","00100000","01100110","00000000","10011100","00000000","00000000","01010110","10010111","01110100","00011111","00000000","00000000","00000000","00000000",
        "00000000","10010101","00000000","00000000","00010001","00000000","00000000","00000000","00000000","10100011","00000000","01100000","00000000","00000000","00000000","00011110",
        "00000000","01101001","10010100","10011010","00000000","01101111","01110011","00000100","10001110","00000000","00000000","10010010","00000000","00000000","00010011","00001101",
        "10000001","00000000","00000000","00000000","00000000","00110111","00000111","00000000","00000000","00000000","10011000","00101000","00000000","00000000","10101011","10000101",
        "00001001","00000000","00011011","00000000","00000000","01000000","00000000","10111011","10100101","00000000","00001100","00111001","00111011","00000000","00000101","00000000",
        "00100111","10101100","00000000","00101111","00000000","10101101","00000000","00111110","10111101","00000000","00000000","00000000","11001101","00000000","00000000","00000000",
        "00010000","00000000","00000000","00101011","00111010","00000000","00000000","00000000","00000000","00100010","00000000","00000000","00000000","00000000","00000000","00000000",
        "01001010","00000000","10111001","01000111","00000000","00000000","00101110","11000000","00000000","00000000","00111000","00000000","01001100","00000000","11010101","00111100",
        "00110100","00000000","00000000","11010010","00000110","00101001","01000101","00110101","00000000","00000000","00000000","11011110","00000000","11100110","00000000","00001000",
        "00000000","00011101","00000000","00000000","00000000","00000000","00000000","00100101","11011100","00000000","00010111","00000000","00011100","00100110","11101010","00011010",
        "00000000","00000011","01000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01101110","01100010","00001110","01110101","00000000",
        "01010001","00000000","00000000","00000000","00000000","00110001","00111101","01010000","00000000","00000000","01011101","00000000","01001111","01010111",
        "01010101","00001011","00010110","00010010","00101100","00000000","00100100","00110110","01011000","00000000","00000000","00000000","01001000","10000000","01101100","00000000",
        "01011111","01110111","00000000","01001011","00000000","00000000","00000000","00011000","10000111","01110010","00000001","01110110","01000011","00000000","00000000","00001010",
        "01100001","00000000","00110011","01001110","00000000","01011001","10001111","00000000","00000000","01011110","00000000","00000000","00000000","01011011","00110000","00000000",
        "00001111","01111100","01001101","01111011","00000010","00000000","01001001","00000000","10000110","00000000","00000000","10011011","00000000","00000000","00010100","00000000",
        "01111101","00000000","00000000","00100000","01100110","00000000","10011100","00000000","00000000","01010110","10010111","01110100","00011111","00000000","00000000","00000000",
        "00000000","00000000","10010101","00000000","00000000","00010001","00000000","00000000","00000000","00000000","10100011","00000000","01100000","00000000","00000000","00000000",
        "00011110","00000000","01101001","10010100","10011010","00000000","01101111","01110011","00000100","10001110","00000000","00000000","10010010","00000000","00000000","00010011",
        "00001101","10000001","00000000","00000000","00000000","00000000","00110111","00000111","00000000","00000000","00000000","10011000","00101000","00000000","00000000","10101011",
        "10000101","00001001","00000000","00011011","00000000","00000000","01000000","00000000","10111011","10100101","00000000","00001100","00111001","00111011","00000000","00000101",
        "00000000","00100111","10101100","00000000","00101111","00000000","10101101","00000000","00111110","10111101","00000000","00000000","00000000","11001101","00000000","00000000",
        "00000000","00010000","00000000","00000000","00101011","00111010","00000000","00000000","00000000","00000000","00100010","00000000","00000000","00000000","00000000","00000000",
        "00000000","01001010","00000000","10111001","01000111","00000000","00000000","00101110","11000000","00000000","00000000","00111000","00000000","01001100","00000000","11010101",
        "00111100","00110100","00000000","00000000","11010010","00000110","00101001","01000101","00110101","00000000","00000000","00000000","11011110","00000000","11100110","00000000",
        "00001000","00000000","00011101","00000000","00000000","00000000","00000000","00000000","00100101","11011100","00000000","00010111","00000000","00011100","00100110","11101010",
        "00011010","00000000","00000011","01000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01101110","01100010","00001110","01110101",
        "00000000","01010001","00000000","00000000","00000000","00000000","00110001","00111101","01010000","00000000","00000000","01011101","00000000","01001111","01010111","01010101",
        "00001011","00010110","00010010","00101100","00000000","00100100","00110110","01011000","00000000","00000000","00000000","01001000","10000000","01101100","00000000","01011111",
        "01110111","00000000","01001011","00000000","00000000","00000000","00011000","10000111","01110010","00000001","01110110","01000011","00000000","00000000","00001010","01100001",
        "00000000","00110011","01001110","00000000","01011001","10001111","00000000","00000000","01011110","00000000","00000000","00000000","01011011","00110000","00000000","00001111",
        "01111100","01001101","01111011","00000010","00000000","01001001","00000000","10000110","00000000","00000000","10011011","00000000","00000000","00010100","00000000","01111101",
        "00000000","00000000","00100000","01100110","00000000","10011100","00000000","00000000","01010110","10010111","01110100","00011111","00000000","00000000","00000000","00000000",
        "00000000","10010101","00000000","00000000","00010001","00000000","00000000","00000000","00000000","10100011","00000000","01100000","00000000","00000000","00000000","00011110",
        "00000000","01101001","10010100","10011010","00000000","01101111","01110011","00000100","10001110","00000000","00000000","10010010","00000000","00000000","00010011","00001101",
        "10000001","00000000","00000000","00000000","00000000","00110111","00000111","00000000","00000000","00000000","10011000","00101000","00000000","00000000","10101011","10000101",
        "00001001","00000000","00011011","00000000","00000000","01000000","00000000","10111011","10100101","00000000","00001100","00111001","00111011","00000000","00000101","00000000",
        "00100111","10101100","00000000","00101111","00000000","10101101","00000000","00111110","10111101","00000000","00000000","00000000","11001101","00000000","00000000","00000000",
        "00010000","00000000","00000000","00101011","00111010","00000000","00000000","00000000","00000000","00100010","00000000","00000000","00000000","00000000","00000000","00000000",
        "01001010","00000000","10111001","01000111","00000000","00000000","00101110","11000000","00000000","00000000","00111000","00000000","01001100","00000000","11010101","00111100",
        "00110100","00000000","00000000","11010010","00000110","00101001","01000101","00110101","00000000","00000000","00000000","11011110","00000000","11100110","00000000","00001000",
        "00000000","00011101","00000000","00000000","00000000","00000000","00000000","00100101","11011100","00000000","00010111","00000000","00011100","00100110","11101010","00011010",
        "00000000","00000011","01000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01101110","01100010","00001110","01110101","00000000",
        "01010001","00000000","00000000","00000000","00000000","00110001","00111101","01010000","00000000","00000000","01011101","00000000","01001111","01010111","01010101",
        "00001011","00010110","00010010","00101100","00000000","00100100","00110110","01011000","00000000","00000000","00000000","01001000","10000000","01101100","00000000","01011111",
        "01110111","00000000","01001011","00000000","00000000","00000000","00011000","10000111","01110010","00000001","01110110","01000011","00000000","00000000","00001010","01100001",
        "00000000","00110011","01001110","00000000","01011001","10001111","00000000","00000000","01011110","00000000","00000000","00000000","01011011","00110000","00000000","00001111",
        "01111100","01001101","01111011","00000010","00000000","01001001","00000000","10000110","00000000","00000000","10011011","00000000","00000000","00010100","00000000","01111101",
        "00000000","00000000","00100000","01100110","00000000","10011100","00000000","00000000","01010110","10010111","01110100","00011111","00000000","00000000","00000000","00000000",
        "00000000","10010101","00000000","00000000","00010001","00000000","00000000","00000000","00000000","10100011","00000000","01100000","00000000","00000000","00000000","00011110",
        "00000000","01101001","10010100","10011010","00000000","01101111","01110011","00000100","10001110","00000000","00000000","10010010","00000000","00000000","00010011","00001101",
        "10000001","00000000","00000000","00000000","00000000","00110111","00000111","00000000","00000000","00000000","10011000","00101000","00000000","00000000","10101011","10000101",
        "00001001","00000000","00011011","00000000","00000000","01000000","00000000","10111011","10100101","00000000","00001100","00111001","00111011","00000000","00000101","00000000",
        "00100111","10101100","00000000","00101111","00000000","10101101","00000000","00111110","10111101","00000000","00000000","00000000","11001101","00000000","00000000","00000000",
        "00010000","00000000","00000000","00101011","00111010","00000000","00000000","00000000","00000000","00100010","00000000","00000000","00000000","00000000","00000000","00000000",
        "01001010","00000000","10111001","01000111","00000000","00000000","00101110","11000000","00000000","00000000","00111000","00000000","01001100","00000000","11010101","00111100",
        "00110100","00000000","00000000","11010010","00000110","00101001","01000101","00110101","00000000","00000000","00000000","11011110","00000000","11100110","00000000","00001000",
        "00000000","00011101","00000000","00000000","00000000","00000000","00000000","00100101","11011100","00000000","00010111","00000000","00011100","00100110","11101010","00011010",
        "00000000","00000011","01000001","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01101110","01100010","00001110","01110101","00000000",
        "01010001","00000000","00000000","00000000","00000000","00110001","00111101","01010000","00000000","00000000","01011101","00000000","01001111","01010111");
constant xxxc_3         : table_4 := (
        "10101010","11110101","11101011","11110000","11010111","00000000","11100001","11010000","10101111","00000000","00000000","00000000","11000011","10001100","10100001","00000000",
        "10110000","10011001","00000000","11000111","00000000","00000000","00000000","11111110","10010000","10100110","00011001","10100100","11011000","00000000","00000000","00010101",
        "10111110","00000000","11101110","11010100","00000000","11001011","10010110","00000000","00000000","11001010","00000000","00000000","00000000","11010001","11111101","00000000",
        "00100001","10110100","11100100","10110111","00110010","00000000","11101100","00000000","10110001","00000000","00000000","10011111","00000000","00000000","00101010","00000000",
        "11000010","00000000","00000000","00100011","11011101","00000000","10101001","00000000","00000000","11110010","10110010","11010110","00101101","00000000","00000000","00000000",
        "00000000","00000000","10111100","00000000","00000000","01000100","00000000","00000000","00000000","00000000","10110110","00000000","11111011","00000000","00000000","00000000",
        "01000010","00000000","11111000","11001110","11001001","00000000","11110110","11110011","01100100","11011010","00000000","00000000","11011001","00000000","00000000","01011100",
        "01100011","11101111","00000000","00000000","00000000","00000000","00111111","01110000","00000000","00000000","00000000","11100010","01010100","00000000","00000000","11010011",
        "11111010","01111000","00000000","01101000","00000000","00000000","01000110","00000000","11001100","11100011","00000000","01111111","01010011","01010010","00000000","10001010",
        "00000000","01101010","11100101","00000000","01100101","00000000","11101000","00000000","01011010","11011011","00000000","00000000","00000000","11001111","00000000","00000000",
        "00000000","10010001","00000000","00000000","01111001","01101011","00000000","00000000","00000000","00000000","10001000","00000000","00000000","00000000","00000000","00000000",
        "00000000","01100111","00000000","11111001","01101101","00000000","00000000","10001001","11110111","00000000","00000000","10000011","00000000","01110001","00000000","11101001",
        "10000100","10001101","00000000","00000000","11110001","10111111","10011101","10000010","10010011","00000000","00000000","00000000","11101101","00000000","11100111","00000000",
        "11001000","00000000","10110101","00000000","00000000","00000000","00000000","00000000","10110011","11111100","00000000","11000100","00000000","11000001","10111000","11110100",
        "11000110","00000000","11011111","10100010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01111110","10001011","11100000","01111010",
        "00000000","10100000","00000000","00000000","00000000","00000000","11000101","10111010","10101000","00000000","00000000","10011110","00000000","10101110","10100111",
        "10101010","11110101","11101011","11110000","11010111","00000000","11100001","11010000","10101111","00000000","00000000","00000000","11000011","10001100","10100001","00000000",
        "10110000","10011001","00000000","11000111","00000000","00000000","00000000","11111110","10010000","10100110","00011001","10100100","11011000","00000000","00000000","00010101",
        "10111110","00000000","11101110","11010100","00000000","11001011","10010110","00000000","00000000","11001010","00000000","00000000","00000000","11010001","11111101","00000000",
        "00100001","10110100","11100100","10110111","00110010","00000000","11101100","00000000","10110001","00000000","00000000","10011111","00000000","00000000","00101010","00000000",
        "11000010","00000000","00000000","00100011","11011101","00000000","10101001","00000000","00000000","11110010","10110010","11010110","00101101","00000000","00000000","00000000",
        "00000000","00000000","10111100","00000000","00000000","01000100","00000000","00000000","00000000","00000000","10110110","00000000","11111011","00000000","00000000","00000000",
        "01000010","00000000","11111000","11001110","11001001","00000000","11110110","11110011","01100100","11011010","00000000","00000000","11011001","00000000","00000000","01011100",
        "01100011","11101111","00000000","00000000","00000000","00000000","00111111","01110000","00000000","00000000","00000000","11100010","01010100","00000000","00000000","11010011",
        "11111010","01111000","00000000","01101000","00000000","00000000","01000110","00000000","11001100","11100011","00000000","01111111","01010011","01010010","00000000","10001010",
        "00000000","01101010","11100101","00000000","01100101","00000000","11101000","00000000","01011010","11011011","00000000","00000000","00000000","11001111","00000000","00000000",
        "00000000","10010001","00000000","00000000","01111001","01101011","00000000","00000000","00000000","00000000","10001000","00000000","00000000","00000000","00000000","00000000",
        "00000000","01100111","00000000","11111001","01101101","00000000","00000000","10001001","11110111","00000000","00000000","10000011","00000000","01110001","00000000","11101001",
        "10000100","10001101","00000000","00000000","11110001","10111111","10011101","10000010","10010011","00000000","00000000","00000000","11101101","00000000","11100111","00000000",
        "11001000","00000000","10110101","00000000","00000000","00000000","00000000","00000000","10110011","11111100","00000000","11000100","00000000","11000001","10111000","11110100",
        "11000110","00000000","11011111","10100010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01111110","10001011","11100000","01111010",
        "00000000","10100000","00000000","00000000","00000000","00000000","11000101","10111010","10101000","00000000","00000000","10011110","00000000","10101110","10100111",
        "10101010","11110101","11101011","11110000","11010111","00000000","11100001","11010000","10101111","00000000","00000000","00000000","11000011","10001100","10100001","00000000",
        "10110000","10011001","00000000","11000111","00000000","00000000","00000000","11111110","10010000","10100110","00011001","10100100","11011000","00000000","00000000","00010101",
        "10111110","00000000","11101110","11010100","00000000","11001011","10010110","00000000","00000000","11001010","00000000","00000000","00000000","11010001","11111101","00000000",
        "00100001","10110100","11100100","10110111","00110010","00000000","11101100","00000000","10110001","00000000","00000000","10011111","00000000","00000000","00101010","00000000",
        "11000010","00000000","00000000","00100011","11011101","00000000","10101001","00000000","00000000","11110010","10110010","11010110","00101101","00000000","00000000","00000000",
        "00000000","00000000","10111100","00000000","00000000","01000100","00000000","00000000","00000000","00000000","10110110","00000000","11111011","00000000","00000000","00000000",
        "01000010","00000000","11111000","11001110","11001001","00000000","11110110","11110011","01100100","11011010","00000000","00000000","11011001","00000000","00000000","01011100",
        "01100011","11101111","00000000","00000000","00000000","00000000","00111111","01110000","00000000","00000000","00000000","11100010","01010100","00000000","00000000","11010011",
        "11111010","01111000","00000000","01101000","00000000","00000000","01000110","00000000","11001100","11100011","00000000","01111111","01010011","01010010","00000000","10001010",
        "00000000","01101010","11100101","00000000","01100101","00000000","11101000","00000000","01011010","11011011","00000000","00000000","00000000","11001111","00000000","00000000",
        "00000000","10010001","00000000","00000000","01111001","01101011","00000000","00000000","00000000","00000000","10001000","00000000","00000000","00000000","00000000","00000000",
        "00000000","01100111","00000000","11111001","01101101","00000000","00000000","10001001","11110111","00000000","00000000","10000011","00000000","01110001","00000000","11101001",
        "10000100","10001101","00000000","00000000","11110001","10111111","10011101","10000010","10010011","00000000","00000000","00000000","11101101","00000000","11100111","00000000",
        "11001000","00000000","10110101","00000000","00000000","00000000","00000000","00000000","10110011","11111100","00000000","11000100","00000000","11000001","10111000","11110100",
        "11000110","00000000","11011111","10100010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01111110","10001011","11100000","01111010",
        "00000000","10100000","00000000","00000000","00000000","00000000","11000101","10111010","10101000","00000000","00000000","10011110","00000000","10101110","10100111",
        "10101010","11110101","11101011","11110000","11010111","00000000","11100001","11010000","10101111","00000000","00000000","00000000","11000011","10001100","10100001","00000000",
        "10110000","10011001","00000000","11000111","00000000","00000000","00000000","11111110","10010000","10100110","00011001","10100100","11011000","00000000","00000000","00010101",
        "10111110","00000000","11101110","11010100","00000000","11001011","10010110","00000000","00000000","11001010","00000000","00000000","00000000","11010001","11111101","00000000",
        "00100001","10110100","11100100","10110111","00110010","00000000","11101100","00000000","10110001","00000000","00000000","10011111","00000000","00000000","00101010","00000000",
        "11000010","00000000","00000000","00100011","11011101","00000000","10101001","00000000","00000000","11110010","10110010","11010110","00101101","00000000","00000000","00000000",
        "00000000","00000000","10111100","00000000","00000000","01000100","00000000","00000000","00000000","00000000","10110110","00000000","11111011","00000000","00000000","00000000",
        "01000010","00000000","11111000","11001110","11001001","00000000","11110110","11110011","01100100","11011010","00000000","00000000","11011001","00000000","00000000","01011100",
        "01100011","11101111","00000000","00000000","00000000","00000000","00111111","01110000","00000000","00000000","00000000","11100010","01010100","00000000","00000000","11010011",
        "11111010","01111000","00000000","01101000","00000000","00000000","01000110","00000000","11001100","11100011","00000000","01111111","01010011","01010010","00000000","10001010",
        "00000000","01101010","11100101","00000000","01100101","00000000","11101000","00000000","01011010","11011011","00000000","00000000","00000000","11001111","00000000","00000000",
        "00000000","10010001","00000000","00000000","01111001","01101011","00000000","00000000","00000000","00000000","10001000","00000000","00000000","00000000","00000000","00000000",
        "00000000","01100111","00000000","11111001","01101101","00000000","00000000","10001001","11110111","00000000","00000000","10000011","00000000","01110001","00000000","11101001",
        "10000100","10001101","00000000","00000000","11110001","10111111","10011101","10000010","10010011","00000000","00000000","00000000","11101101","00000000","11100111","00000000",
        "11001000","00000000","10110101","00000000","00000000","00000000","00000000","00000000","10110011","11111100","00000000","11000100","00000000","11000001","10111000","11110100",
        "11000110","00000000","11011111","10100010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01111110","10001011","11100000","01111010",
        "00000000","10100000","00000000","00000000","00000000","00000000","11000101","10111010","10101000","00000000","00000000","10011110","00000000","10101110","10100111",
        "10101010","11110101","11101011","11110000","11010111","00000000","11100001","11010000","10101111","00000000","00000000","00000000","11000011","10001100","10100001","00000000",
        "10110000","10011001","00000000","11000111","00000000","00000000","00000000","11111110","10010000","10100110","00011001","10100100","11011000","00000000","00000000","00010101",
        "10111110","00000000","11101110","11010100","00000000","11001011","10010110","00000000","00000000","11001010","00000000","00000000","00000000","11010001","11111101","00000000",
        "00100001","10110100","11100100","10110111","00110010","00000000","11101100","00000000","10110001","00000000","00000000","10011111","00000000","00000000","00101010","00000000",
        "11000010","00000000","00000000","00100011","11011101","00000000","10101001","00000000","00000000","11110010","10110010","11010110","00101101","00000000","00000000","00000000",
        "00000000","00000000","10111100","00000000","00000000","01000100","00000000","00000000","00000000","00000000","10110110","00000000","11111011","00000000","00000000","00000000",
        "01000010","00000000","11111000","11001110","11001001","00000000","11110110","11110011","01100100","11011010","00000000","00000000","11011001","00000000","00000000","01011100",
        "01100011","11101111","00000000","00000000","00000000","00000000","00111111","01110000","00000000","00000000","00000000","11100010","01010100","00000000","00000000","11010011",
        "11111010","01111000","00000000","01101000","00000000","00000000","01000110","00000000","11001100","11100011","00000000","01111111","01010011","01010010","00000000","10001010",
        "00000000","01101010","11100101","00000000","01100101","00000000","11101000","00000000","01011010","11011011","00000000","00000000","00000000","11001111","00000000","00000000",
        "00000000","10010001","00000000","00000000","01111001","01101011","00000000","00000000","00000000","00000000","10001000","00000000","00000000","00000000","00000000","00000000",
        "00000000","01100111","00000000","11111001","01101101","00000000","00000000","10001001","11110111","00000000","00000000","10000011","00000000","01110001","00000000","11101001",
        "10000100","10001101","00000000","00000000","11110001","10111111","10011101","10000010","10010011","00000000","00000000","00000000","11101101","00000000","11100111","00000000",
        "11001000","00000000","10110101","00000000","00000000","00000000","00000000","00000000","10110011","11111100","00000000","11000100","00000000","11000001","10111000","11110100",
        "11000110","00000000","11011111","10100010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01111110","10001011","11100000","01111010",
        "00000000","10100000","00000000","00000000","00000000","00000000","11000101","10111010","10101000","00000000","00000000","10011110","00000000","10101110","10100111",
        "10101010","11110101","11101011","11110000","11010111","00000000","11100001","11010000","10101111","00000000","00000000","00000000","11000011","10001100","10100001","00000000",
        "10110000","10011001","00000000","11000111","00000000","00000000","00000000","11111110","10010000","10100110","00011001","10100100","11011000","00000000","00000000","00010101",
        "10111110","00000000","11101110","11010100","00000000","11001011","10010110","00000000","00000000","11001010","00000000","00000000","00000000","11010001","11111101","00000000",
        "00100001","10110100","11100100","10110111","00110010","00000000","11101100","00000000","10110001","00000000","00000000","10011111","00000000","00000000","00101010","00000000",
        "11000010","00000000","00000000","00100011","11011101","00000000","10101001","00000000","00000000","11110010","10110010","11010110","00101101","00000000","00000000","00000000",
        "00000000","00000000","10111100","00000000","00000000","01000100","00000000","00000000","00000000","00000000","10110110","00000000","11111011","00000000","00000000","00000000",
        "01000010","00000000","11111000","11001110","11001001","00000000","11110110","11110011","01100100","11011010","00000000","00000000","11011001","00000000","00000000","01011100",
        "01100011","11101111","00000000","00000000","00000000","00000000","00111111","01110000","00000000","00000000","00000000","11100010","01010100","00000000","00000000","11010011",
        "11111010","01111000","00000000","01101000","00000000","00000000","01000110","00000000","11001100","11100011","00000000","01111111","01010011","01010010","00000000","10001010",
        "00000000","01101010","11100101","00000000","01100101","00000000","11101000","00000000","01011010","11011011","00000000","00000000","00000000","11001111","00000000","00000000",
        "00000000","10010001","00000000","00000000","01111001","01101011","00000000","00000000","00000000","00000000","10001000","00000000","00000000","00000000","00000000","00000000",
        "00000000","01100111","00000000","11111001","01101101","00000000","00000000","10001001","11110111","00000000","00000000","10000011","00000000","01110001","00000000","11101001",
        "10000100","10001101","00000000","00000000","11110001","10111111","10011101","10000010","10010011","00000000","00000000","00000000","11101101","00000000","11100111","00000000",
        "11001000","00000000","10110101","00000000","00000000","00000000","00000000","00000000","10110011","11111100","00000000","11000100","00000000","11000001","10111000","11110100",
        "11000110","00000000","11011111","10100010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01111110","10001011","11100000","01111010",
        "00000000","10100000","00000000","00000000","00000000","00000000","11000101","10111010","10101000","00000000","00000000","10011110","00000000","10101110","10100111",
        "10101010","11110101","11101011","11110000","11010111","00000000","11100001","11010000","10101111","00000000","00000000","00000000","11000011","10001100","10100001","00000000",
        "10110000","10011001","00000000","11000111","00000000","00000000","00000000","11111110","10010000","10100110","00011001","10100100","11011000","00000000","00000000","00010101",
        "10111110","00000000","11101110","11010100","00000000","11001011","10010110","00000000","00000000","11001010","00000000","00000000","00000000","11010001","11111101","00000000",
        "00100001","10110100","11100100","10110111","00110010","00000000","11101100","00000000","10110001","00000000","00000000","10011111","00000000","00000000","00101010","00000000",
        "11000010","00000000","00000000","00100011","11011101","00000000","10101001","00000000","00000000","11110010","10110010","11010110","00101101","00000000","00000000","00000000",
        "00000000","00000000","10111100","00000000","00000000","01000100","00000000","00000000","00000000","00000000","10110110","00000000","11111011","00000000","00000000","00000000",
        "01000010","00000000","11111000","11001110","11001001","00000000","11110110","11110011","01100100","11011010","00000000","00000000","11011001","00000000","00000000","01011100",
        "01100011","11101111","00000000","00000000","00000000","00000000","00111111","01110000","00000000","00000000","00000000","11100010","01010100","00000000","00000000","11010011",
        "11111010","01111000","00000000","01101000","00000000","00000000","01000110","00000000","11001100","11100011","00000000","01111111","01010011","01010010","00000000","10001010",
        "00000000","01101010","11100101","00000000","01100101","00000000","11101000","00000000","01011010","11011011","00000000","00000000","00000000","11001111","00000000","00000000",
        "00000000","10010001","00000000","00000000","01111001","01101011","00000000","00000000","00000000","00000000","10001000","00000000","00000000","00000000","00000000","00000000",
        "00000000","01100111","00000000","11111001","01101101","00000000","00000000","10001001","11110111","00000000","00000000","10000011","00000000","01110001","00000000","11101001",
        "10000100","10001101","00000000","00000000","11110001","10111111","10011101","10000010","10010011","00000000","00000000","00000000","11101101","00000000","11100111","00000000",
        "11001000","00000000","10110101","00000000","00000000","00000000","00000000","00000000","10110011","11111100","00000000","11000100","00000000","11000001","10111000","11110100",
        "11000110","00000000","11011111","10100010","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","01111110","10001011","11100000","01111010",
        "00000000","10100000","00000000","00000000","00000000","00000000","11000101","10111010","10101000","00000000","00000000","10011110","00000000","10101110","10100111");
------------------------------------------------------------------------------------------------------------
--CLK 0
signal s1_in             : std_logic_vector(7 downto 0);
signal s3_in             : std_logic_vector(7 downto 0);
signal hard_input_in     : std_logic_vector(255 downto 0);
signal soft_input_in     : input_data_array(255 downto 0);
------------------------------------------------------------------------------------------------------------
--CLK 1
type state_machine is (no_error_state, one_error_state, two_error_state, unable_to_correct_state);
signal state    	 : state_machine := unable_to_correct_state;
signal s1_temp           : std_logic_vector(7 downto 0); -- maximum 255
signal s3_temp           : std_logic_vector(7 downto 0);
signal s1_flag           : std_logic; 
signal s3_flag           : std_logic;
signal hard_input_pass_1 : std_logic_vector(255 downto 0);
signal soft_input_1      : input_data_array(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 2
signal soft_input_2      : input_data_array(255 downto 0);
signal s1_temp_1         : std_logic_vector(7 downto 0);
signal s3_temp_1         : std_logic_vector(7 downto 0);
signal s1_flag_1         : std_logic; 
signal s3_flag_1         : std_logic;
signal s1_plus_1         : std_logic_vector(7 downto 0);
signal sum_1_1           : std_logic_vector(8 downto 0);
signal sum_1_2           : std_logic_vector(8 downto 0);
signal sum_1_3           : std_logic_vector(8 downto 0);
signal sum_1_4           : std_logic_vector(8 downto 0); -- Maximum 256
signal hard_input_pass_2 : std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 3
signal soft_input_3     : input_data_array(255 downto 0);
signal s1_plus_1_pass1  : std_logic_vector(7 downto 0);
signal log_s1_plus_1    : std_logic_vector(8 downto 0);
signal s3_temp_2        : std_logic_vector(7 downto 0);
signal s1_temp_2        : std_logic_vector(7 downto 0);
signal s1_s3_flag       : std_logic;
signal sum_2_1          : std_logic_vector(8 downto 0);
signal sum_2_2          : std_logic_vector(8 downto 0);
signal sum_2_3          : std_logic_vector(8 downto 0);
signal sum_2_4          : std_logic_vector(8 downto 0);
signal sum_2_5          : std_logic_vector(8 downto 0);
signal hard_input_pass_3: std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 4
signal soft_input_4     : input_data_array(255 downto 0);
signal s1_plus_1_pass2  : std_logic_vector(7 downto 0);
signal log_s1_plus_1m2  : std_logic_vector(8 downto 0); -- because of shifting, just in case
signal log_s1_plus_2    : std_logic_vector(8 downto 0);
signal s3_temp_3        : std_logic_vector(7 downto 0);
signal s1_temp_3        : std_logic_vector(7 downto 0);
signal s1_s3_flag_1     : std_logic;
signal sum_3_1          : std_logic_vector(8 downto 0);
signal sum_3_2          : std_logic_vector(8 downto 0);
signal sum_3_3          : std_logic_vector(8 downto 0);
signal sum_3_4          : std_logic_vector(8 downto 0);
signal sum_3_5          : std_logic_vector(8 downto 0);
signal hard_input_pass_4: std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 5
signal soft_input_5        : input_data_array(255 downto 0);
signal s1_plus_1_pass3     : std_logic_vector(7 downto 0);
signal s1_power3_log       : std_logic_vector(9 downto 0); -- because of adding, just in case  
signal log_s1_plus_1m2_exp : std_logic_vector(9 downto 0);
signal log_s1_plus_2_exp   : std_logic_vector(9 downto 0); 
signal s3_temp_4           : std_logic_vector(7 downto 0);
signal s1_temp_4           : std_logic_vector(7 downto 0);
signal s1_s3_flag_2        : std_logic;
signal sum_4_1             : std_logic_vector(8 downto 0);
signal sum_4_2             : std_logic_vector(8 downto 0);
signal sum_4_3             : std_logic_vector(8 downto 0);
signal sum_4_4             : std_logic_vector(8 downto 0);
signal sum_4_5             : std_logic_vector(8 downto 0);
signal hard_input_pass_5   : std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 6
signal soft_input_6     : input_data_array(255 downto 0);
signal s1_plus_1_pass4  : std_logic_vector(7 downto 0); 
signal s1_power3_temp   : std_logic_vector(7 downto 0); -- temp value of s1_power3, after adding 1 it will be complete
signal s3_temp_5        : std_logic_vector(7 downto 0);       
signal s1_temp_5        : std_logic_vector(7 downto 0);       
signal s1_s3_flag_3     : std_logic;     
signal s1_power3_log_1  : std_logic_vector(9 downto 0);
signal sum_5_1          : std_logic_vector(8 downto 0);
signal sum_5_2          : std_logic_vector(8 downto 0);
signal sum_5_3          : std_logic_vector(8 downto 0);
signal sum_5_4          : std_logic_vector(8 downto 0);
signal sum_5_5          : std_logic_vector(8 downto 0);
signal hard_input_pass_6: std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 7
signal soft_input_7     : input_data_array(255 downto 0);
signal s1_plus_1_pass5  : std_logic_vector(7 downto 0);
signal s1_power3        : std_logic_vector(7 downto 0); -- only adding 1, no need to change
signal s1_power3_log_2  : std_logic_vector(9 downto 0);
signal s3_temp_6        : std_logic_vector(7 downto 0); 
signal s1_temp_6        : std_logic_vector(7 downto 0); 
signal s1_s3_flag_4     : std_logic;   
signal sum_6_1          : std_logic_vector(8 downto 0);
signal sum_6_2          : std_logic_vector(8 downto 0);
signal sum_6_3          : std_logic_vector(8 downto 0);
signal sum_6_4          : std_logic_vector(8 downto 0);
signal sum_6_5          : std_logic_vector(8 downto 0);
signal hard_input_pass_7: std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 8
signal soft_input_8     : input_data_array(255 downto 0);
signal s1_plus_1_pass6  : std_logic_vector(7 downto 0);
signal s1_power3_1      : std_logic_vector(7 downto 0);
signal s1_power3_log_3  : std_logic_vector(9 downto 0);
signal s3_temp_7        : std_logic_vector(7 downto 0);
signal s1_temp_7        : std_logic_vector(7 downto 0);
signal A_index          : std_logic_vector(8 downto 0); -- s1_power3 xor s3_temp_6, but maybe 9 bits is enough
signal s1_s3_flag_5     : std_logic; 
signal s1_power3_s3_flag: std_logic; 
signal s1_power3_exp    : std_logic_vector(8 downto 0);
signal s3_temp_6_exp    : std_logic_vector(8 downto 0);
signal sum_7_1          : std_logic_vector(8 downto 0);
signal sum_7_2          : std_logic_vector(8 downto 0);
signal sum_7_3          : std_logic_vector(8 downto 0);
signal sum_7_4          : std_logic_vector(8 downto 0);
signal sum_7_5          : std_logic_vector(8 downto 0);
signal hard_input_pass_8: std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 9
signal soft_input_9       : input_data_array(255 downto 0);
signal s1_plus_1_pass7    : std_logic_vector(7 downto 0);
signal s1_power3_2        : std_logic_vector(7 downto 0);
signal s3_temp_8          : std_logic_vector(7 downto 0);
signal s1_temp_8          : std_logic_vector(7 downto 0);
signal A                  : std_logic_vector(9 downto 0); -- up to 1024, should be enough
signal s1_s3_flag_6       : std_logic; 
signal s1_power3_s3_flag_1: std_logic; 
signal sum_8_1            : std_logic_vector(8 downto 0);
signal sum_8_2            : std_logic_vector(8 downto 0);
signal sum_8_3            : std_logic_vector(8 downto 0);
signal sum_8_4            : std_logic_vector(8 downto 0);
signal sum_8_5            : std_logic_vector(8 downto 0);
signal hard_input_pass_9  : std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 10
signal soft_input_10      : input_data_array(255 downto 0);
signal s1_plus_1_pass8    : std_logic_vector(7 downto 0);
signal s1_power3_3        : std_logic_vector(7 downto 0);
signal s3_temp_9          : std_logic_vector(7 downto 0);
signal s1_temp_9          : std_logic_vector(7 downto 0);
signal xxxc1a             : std_logic_vector(1 downto 0);
signal xxxc2a             : std_logic_vector(7 downto 0);
signal xxxc3a             : std_logic_vector(7 downto 0);
signal s1_s3_flag_7       : std_logic; 
signal s1_power3_s3_flag_2: std_logic; 
signal log_v              : std_logic_vector(8 downto 0);
signal s1_power3_log_4    : std_logic_vector(9 downto 0); 
signal sum_9_1            : std_logic_vector(8 downto 0);
signal sum_9_2            : std_logic_vector(8 downto 0);
signal sum_9_3            : std_logic_vector(8 downto 0);
signal sum_9_4            : std_logic_vector(8 downto 0);
signal sum_9_5            : std_logic_vector(8 downto 0);
signal hard_input_pass_10 : std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 11
signal soft_input_11      : input_data_array(255 downto 0);
signal s1_plus_1_pass9    : std_logic_vector(7 downto 0);
signal s1_power3_4        : std_logic_vector(7 downto 0);
signal s3_temp_10         : std_logic_vector(7 downto 0);
signal s1_temp_10         : std_logic_vector(7 downto 0);
signal flag_1             : std_logic; 
signal flag_2             : std_logic; 
signal xxxc2a_1           : std_logic_vector(7 downto 0);
signal xxxc3a_1           : std_logic_vector(7 downto 0);
signal s1_s3_flag_8       : std_logic; 
signal s1_power3_s3_flag_3: std_logic; 
signal log_table_value_s1p: std_logic_vector(8 downto 0);
signal A_temp             : integer;
signal sum_10_1           : std_logic_vector(8 downto 0);
signal sum_10_2           : std_logic_vector(8 downto 0);
signal sum_10_3           : std_logic_vector(8 downto 0);
signal sum_10_4           : std_logic_vector(8 downto 0);
signal sum_10_5           : std_logic_vector(8 downto 0);
signal hard_input_pass_11 : std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 12
signal soft_input_12      : input_data_array(255 downto 0);
signal s1_plus_1_pass10   : std_logic_vector(7 downto 0);
signal eh1_temp           : integer;
signal eh2_temp           : integer;
signal eh3_temp           : integer;
signal s3_temp_11         : std_logic_vector(7 downto 0);
signal s1_temp_11         : std_logic_vector(7 downto 0);
signal s1_s3_flag_9       : std_logic;  
signal sum_11_1           : std_logic_vector(8 downto 0);
signal sum_11_2           : std_logic_vector(8 downto 0);
signal sum_11_3           : std_logic_vector(8 downto 0);
signal sum_11_4           : std_logic_vector(8 downto 0);
signal sum_11_5           : std_logic_vector(8 downto 0);
signal hard_input_pass_12 : std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 13
signal soft_input_13      : input_data_array(255 downto 0);
signal s1_plus_1_pass11   : std_logic_vector(7 downto 0);
signal s3_temp_12         : std_logic_vector(7 downto 0);
signal s1_temp_12         : std_logic_vector(7 downto 0);
signal s1_s3_flag_10      : std_logic;
signal s1_power3_5        : std_logic_vector(7 downto 0);
signal s1_power3_s3_flag_4: std_logic;
signal sum_12_1           : std_logic_vector(8 downto 0);
signal sum_12_2           : std_logic_vector(8 downto 0);
signal sum_12_3           : std_logic_vector(8 downto 0);
signal sum_12_4           : std_logic_vector(8 downto 0);
signal sum_12_5           : std_logic_vector(8 downto 0);
signal hard_input_pass_13 : std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 14
signal soft_input_14        : input_data_array(255 downto 0);
signal s3_temp_13           : std_logic_vector(7 downto 0);
signal s1_temp_13           : std_logic_vector(7 downto 0);
signal s1_power3_6          : std_logic_vector(7 downto 0);
signal s1_s3_flag_11        : std_logic;
signal s1_power3_s3_flag_5  : std_logic; 
signal indi_1               : boolean; 
signal indi_2               : boolean; 
signal sum_13_1             : std_logic_vector(8 downto 0);
signal sum_13_2             : std_logic_vector(8 downto 0);
signal sum_13_3             : std_logic_vector(8 downto 0);
signal sum_13_4             : std_logic_vector(8 downto 0);
signal sum_13_5             : std_logic_vector(8 downto 0);
signal hard_input_pass_14   : std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 15
signal soft_input_15         : input_data_array(255 downto 0);
signal log_table_value_s1p_1 : std_logic_vector(8 downto 0);
signal s1_power3_7           : std_logic_vector(7 downto 0);
signal s3_temp_14            : std_logic_vector(7 downto 0);
signal xxxc2a_2              : std_logic_vector(7 downto 0);
signal xxxc3a_2              : std_logic_vector(7 downto 0);
signal s1_s3_flag_12         : std_logic; 
signal s1_power3_s3_flag_6   : std_logic; 
signal sum_14_1              : std_logic_vector(8 downto 0);
signal sum_14_2              : std_logic_vector(8 downto 0);
signal sum_14_3              : std_logic_vector(8 downto 0);
signal sum_14_4              : std_logic_vector(8 downto 0);
signal sum_14_5              : std_logic_vector(8 downto 0);
signal hard_input_pass_15    : std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 16
signal soft_input_16         : input_data_array(255 downto 0);
signal sum_15_1              : std_logic_vector(8 downto 0);
signal sum_15_2              : std_logic_vector(8 downto 0);
signal sum_15_3              : std_logic_vector(8 downto 0);
signal sum_15_4              : std_logic_vector(8 downto 0);
signal sum_15_5              : std_logic_vector(8 downto 0);
signal hard_input_pass_16    : std_logic_vector(255 downto 0);
-------------------------------------------------------------------------------------------------------------
--CLK 17
signal soft_input_17         : input_data_array(255 downto 0);
signal hard_input_f          : std_logic_vector(255 downto 0);  
signal next_state            : state_machine;
signal eh1_n1                : integer;
signal eh1_n2                : integer;
signal eh1                   : integer;   
signal eh2                   : integer;               
signal eh3                   : integer;     
signal sum_16_1              : std_logic_vector(8 downto 0);
signal sum_16_2              : std_logic_vector(8 downto 0);
signal sum_16_3              : std_logic_vector(8 downto 0);
signal sum_16_4              : std_logic_vector(8 downto 0);
signal sum_16_5              : std_logic_vector(8 downto 0);     
-------------------------------------------------------------------------------------------------------------
--CLK 18
signal soft_input_18         : input_data_array(255 downto 0);
signal next_state_1          : state_machine;
signal hard_output_temp      : std_logic_vector(255 downto 0);  
signal eh1_pass              : integer;            
signal eh2_pass              : integer;      
signal eh3_pass              : integer;             
signal eh1_pass_n1           : integer;      
signal eh1_pass_n2           : integer;      
signal eh2_pass_n1           : integer;      
signal eh3_pass_n1           : integer;      
signal sum_16_temp_1         : std_logic_vector(8 downto 0);              
-------------------------------------------------------------------------------------------------------------
--CLK 19     
signal soft_input_19           : input_data_array(255 downto 0);  
signal next_state_2            : state_machine;  
signal hard_output_error_1     : std_logic; 
signal hard_output_error_2     : std_logic; 
signal hard_output_error_3     : std_logic; 
signal hard_output_error_rest_1: std_logic_vector(255 downto 0);  
signal eh1_pass_1              : integer;
signal eh2_pass_1              : integer;
signal eh3_pass_1              : integer;
signal eh2_pass_n2_1           : integer;
signal eh3_pass_n2_1           : integer;
signal eh1_pass_n1_1           : integer;
signal eh2_pass_n1_1           : integer;
signal eh3_pass_n1_1           : integer;
-------------------------------------------------------------------------------------------------------------
--CLK 20
signal soft_input_20           : input_data_array(255 downto 0);
signal hard_output_error_rest_2: std_logic_vector(255 downto 0);  
signal error_position_temp     : output_error_location_array(2 downto 0); 
signal corrections_temp        : std_logic_vector(2 downto 0); 
-------------------------------------------------------------------------------------------------------------
--CLK 21
signal soft_input_21           : input_data_array(255 downto 0);
signal indi_3                  : boolean;
signal hard_output_error_rest_3: std_logic_vector(255 downto 0);  
signal last_bit                : std_logic;      
signal error_position_temp_1   : output_error_location_array(2 downto 0); 
signal corrections_temp_1      : std_logic_vector(2 downto 0);        
-------------------------------------------------------------------------------------------------------------
--CLK 22
signal soft_input_22           : input_data_array(255 downto 0);
signal indi_4                  : boolean;
signal hard_output_error_rest_4: std_logic_vector(255 downto 0);  
signal last_bit_1              : std_logic;      
signal error_position_temp_2   : output_error_location_array(2 downto 0); 
signal corrections_temp_2      : std_logic_vector(2 downto 0);      
-------------------------------------------------------------------------------------------------------------
--CLK 23
signal soft_input_23           : input_data_array(255 downto 0);
signal hard_output_error_rest_5: std_logic_vector(255 downto 0);  
signal error_position_temp_3   : output_error_location_array(2 downto 0);
signal corrections_temp_3      : std_logic_vector(2 downto 0);         
-------------------------------------------------------------------------------------------------------------
--CLK 24
signal soft_input_24           : input_data_array(255 downto 0);
signal hard_output_error_rest_6: std_logic_vector(255 downto 0); 
signal error_position_temp_4   : output_error_location_array(2 downto 0); 
signal corrections_temp_4      : std_logic_vector(2 downto 0);    
-------------------------------------------------------------------------------------------------------------
--CLK 25
signal soft_input_25           : input_data_array(255 downto 0);
signal hard_output_error_rest_7: std_logic_vector(255 downto 0); 
signal error_position_temp_5   : output_error_location_array(2 downto 0); 
signal corrections_temp_5      : std_logic_vector(2 downto 0);   
-------------------------------------------------------------------------------------------------------------
--CLK 26
signal soft_input_26           : input_data_array(255 downto 0);
signal hard_output_error_rest_8: std_logic_vector(255 downto 0); 
signal error_position_temp_6   : output_error_location_array(2 downto 0); 
signal corrections_temp_6      : std_logic_vector(2 downto 0);   
-------------------------------------------------------------------------------------------------------------
--CLK 27
signal soft_input_27           : input_data_array(255 downto 0);
signal hard_output_error_rest_9: std_logic_vector(255 downto 0); 
signal error_position_temp_7   : output_error_location_array(2 downto 0); 
signal corrections_temp_7      : std_logic_vector(2 downto 0);   
-------------------------------------------------------------------------------------------------------------
--CLK 28
signal soft_input_28            : input_data_array(255 downto 0);
signal hard_output_error_rest_10: std_logic_vector(255 downto 0); 
signal error_position_temp_8    : output_error_location_array(2 downto 0); 
signal corrections_temp_8       : std_logic_vector(2 downto 0);   
-------------------------------------------------------------------------------------------------------------
--CLK 29
signal soft_input_29            : input_data_array(255 downto 0);
signal hard_output_error_rest_11: std_logic_vector(255 downto 0); 
signal error_position_temp_9    : output_error_location_array(2 downto 0); 
signal corrections_temp_9       : std_logic_vector(2 downto 0);   
-------------------------------------------------------------------------------------------------------------
--CLK 30
signal soft_input_30            : input_data_array(255 downto 0);
signal hard_output_error_rest_12: std_logic_vector(255 downto 0); 
signal error_position_temp_10   : output_error_location_array(2 downto 0); 
signal corrections_temp_10      : std_logic_vector(2 downto 0); 
-------------------------------------------------------------------------------------------------------------
--CLK 31
signal soft_input_31            : input_data_array(255 downto 0);
signal hard_output_error_rest_13: std_logic_vector(255 downto 0); 
signal error_position_temp_11   : output_error_location_array(2 downto 0); 
signal corrections_temp_11      : std_logic_vector(2 downto 0); 
-------------------------------------------------------------------------------------------------------------
--CLK 32
signal soft_input_32            : input_data_array(255 downto 0);
signal hard_output_error_rest_14: std_logic_vector(255 downto 0); 
signal error_position_temp_12   : output_error_location_array(2 downto 0); 
signal corrections_temp_12      : std_logic_vector(2 downto 0); 
-------------------------------------------------------------------------------------------------------------
--CLK 33
signal soft_input_33            : input_data_array(255 downto 0);
signal hard_output_error_rest_15: std_logic_vector(255 downto 0); 
signal error_position_temp_13   : output_error_location_array(2 downto 0); 
signal corrections_temp_13      : std_logic_vector(2 downto 0); 
-------------------------------------------------------------------------------------------------------------
--CLK 34
signal soft_input_34            : input_data_array(255 downto 0);
signal hard_output_error_rest_16: std_logic_vector(255 downto 0); 
signal error_position_temp_14   : output_error_location_array(2 downto 0); 
signal corrections_temp_14      : std_logic_vector(2 downto 0); 
-------------------------------------------------------------------------------------------------------------
--CLK 35
signal soft_input_35            : input_data_array(255 downto 0);
signal hard_output_error_rest_17: std_logic_vector(255 downto 0); 
signal error_position_temp_15   : output_error_location_array(2 downto 0); 
signal corrections_temp_15      : std_logic_vector(2 downto 0); 
-------------------------------------------------------------------------------------------------------------
--CLK 36
signal soft_input_36            : input_data_array(255 downto 0);
signal hard_output_error_rest_18: std_logic_vector(255 downto 0); 
signal error_position_temp_16   : output_error_location_array(2 downto 0); 
signal corrections_temp_16      : std_logic_vector(2 downto 0); 
-------------------------------------------------------------------------------------------------------------
--CLK 37
signal soft_input_37            : input_data_array(255 downto 0);
signal hard_output_error_rest_19: std_logic_vector(255 downto 0); 
signal error_position_temp_17   : output_error_location_array(2 downto 0); 
signal corrections_temp_17      : std_logic_vector(2 downto 0); 
-------------------------------------------------------------------------------------------------------------
--CLK 38
signal soft_input_38            : input_data_array(255 downto 0);
signal hard_output_error_rest_20: std_logic_vector(255 downto 0); 
signal error_position_temp_18   : output_error_location_array(2 downto 0); 
signal corrections_temp_18      : std_logic_vector(2 downto 0); 
-------------------------------------------------------------------------------------------------------------
--CLK 39
signal soft_input_39            : input_data_array(255 downto 0);
signal hard_output_error_rest_21: std_logic_vector(255 downto 0); 
signal error_position_temp_19   : output_error_location_array(2 downto 0); 
signal corrections_temp_19      : std_logic_vector(2 downto 0); 
-------------------------------------------------------------------------------------------------------------
--CLK 40
signal soft_input_40            : input_data_array(255 downto 0);
signal hard_output_error_rest_22: std_logic_vector(255 downto 0); 
signal error_position_temp_20   : output_error_location_array(2 downto 0); 
signal corrections_temp_20      : std_logic_vector(2 downto 0); 

begin
------------------------------------------------------------------------------------------------------------
-- Define processes : (CLK 0)
------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                soft_input_in        <= (others => (others => '0'));
                hard_input_in        <= (others => '0');
                s1_in                <= (others => '0');
                s3_in                <= (others => '0');
        elsif rising_edge(clk) then
                soft_input_in        <= soft_input;
                hard_input_in        <= hard_input;
                s1_in                <= s1;
                s3_in                <= s3;
        end if;
end process;
------------------------------------------------------------------------------------------------------------
-- Define processes : Get data into the design (CLK 1)
------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_temp           <= (others => '0');
                s3_temp           <= (others => '0');
                s1_flag           <= '0';
                s3_flag           <= '0';
                hard_input_pass_1 <= (others => '0');
                soft_input_1      <= (others => (others => '0'));
        elsif rising_edge(clk) then
                soft_input_1      <= soft_input_in;
                hard_input_pass_1 <= hard_input_in;
                s1_temp           <= s1_in; -- Store the first s1 and s3
                s3_temp           <= s3_in;
                if (s1_in = "00000000") then
                        s1_flag <= '1';
                else
                        s1_flag <= '0';
                end if;
                if (s3_in = "00000000") then
                        s3_flag <= '1';
                else
                        s3_flag <= '0';
                end if;
        end if;
end process;
------------------------------------------------------------------------------------------------------------
-- Define processes : (CLK 2)
------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1   	 <= "00000001"; 
                s3_temp_1        <= (others => '0');
                s1_temp_1        <= (others => '0');
                s1_flag_1        <= '0';
                s3_flag_1        <= '0';
                hard_input_pass_2<= (others => '0'); 
                soft_input_2     <= (others => (others => '0'));
        elsif rising_edge(clk) then   
                soft_input_2     <= soft_input_1;      
                hard_input_pass_2<= hard_input_pass_1;
                s1_plus_1   	 <= s1_temp;
                s3_temp_1        <= s3_temp;     -- s3 
                s1_temp_1        <= s1_temp;     -- s1 
                s1_flag_1        <= s1_flag;
                s3_flag_1        <= s3_flag;
        end if;
end process;
------------------------------------------------------------------------------------------------------------
-- Define processes : (CLK 3)
------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1_pass1   <= (others => '0');
                log_s1_plus_1     <= "000000001";
                s3_temp_2         <= (others => '0');
                s1_temp_2         <= (others => '0');
                s1_s3_flag        <= '0';
                hard_input_pass_3 <= (others => '0'); 
                soft_input_3      <= (others => (others => '0'));
        elsif rising_edge(clk) then  
                soft_input_3      <= soft_input_2;  
                hard_input_pass_3 <= hard_input_pass_2;
                s1_plus_1_pass1   <= s1_plus_1;
                log_s1_plus_1     <= log_table(to_integer(unsigned(s1_plus_1)));
                s3_temp_2         <= s3_temp_1;
                s1_temp_2         <= s1_temp_1;
                s1_s3_flag        <= s1_flag_1 and s3_flag_1; -- s1 == s3 = 0, no error
        end if;
end process;
------------------------------------------------------------------------------------------------------------
-- Define processes : (CLK 4)
------------------------------------------------------------------------------------------------------------
--process(clk, reset, start)
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1_pass2  <= (others => '0');
                log_s1_plus_2    <= (others => '0');
                log_s1_plus_1m2  <= (others => '0');
                s3_temp_3        <= (others => '0');
                s1_temp_3        <= (others => '0');
                s1_s3_flag_1     <= '0';
                hard_input_pass_4<= (others => '0'); 
                soft_input_4     <= (others => (others => '0'));
        elsif rising_edge(clk) then  
                soft_input_4     <= soft_input_3;  
                hard_input_pass_4<= hard_input_pass_3;
                s1_plus_1_pass2  <= s1_plus_1_pass1;
                log_s1_plus_1m2  <= std_logic_vector(shift_left(unsigned(log_s1_plus_1), 1));
                log_s1_plus_2    <= log_s1_plus_1;
                s3_temp_3        <= s3_temp_2;
                s1_temp_3        <= s1_temp_2;
                s1_s3_flag_1     <= s1_s3_flag;
        end if;
end process;
------------------------------------------------------------------------------------------------------------
-- Define processes : (CLK 5)
------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1_pass3        <= (others => '0');
                log_s1_plus_1m2_exp    <= (others => '0');
                log_s1_plus_2_exp      <= (others => '0');
                s3_temp_4              <= (others => '0');
                s1_temp_4              <= (others => '0');
                s1_s3_flag_2           <= '0';
                hard_input_pass_5      <= (others => '0'); 
                soft_input_5           <= (others => (others => '0'));
        elsif rising_edge(clk) then  
                soft_input_5           <= soft_input_4;
                hard_input_pass_5      <= hard_input_pass_4;
                s1_plus_1_pass3        <= s1_plus_1_pass2;
                log_s1_plus_1m2_exp    <= ('0' & log_s1_plus_1m2);
                log_s1_plus_2_exp      <= ('0' & log_s1_plus_2); 
                s3_temp_4              <= s3_temp_3;
                s1_temp_4              <= s1_temp_3;
                s1_s3_flag_2           <= s1_s3_flag_1;
        end if;
end process;
------------------------------------------------------------------------------------------------------------
-- Define processes : (CLK 6)
------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1_pass4        <= "00000001";
                s1_power3_log          <= "0000000001";
                s3_temp_5              <= (others => '0');
                s1_temp_5              <= (others => '0');
                s1_s3_flag_3           <= '0';
                hard_input_pass_6      <= (others => '0');
                soft_input_6           <= (others => (others => '0')); 
        elsif rising_edge(clk) then  
                soft_input_6           <= soft_input_5;
                hard_input_pass_6      <= hard_input_pass_5;
                s1_plus_1_pass4        <= s1_plus_1_pass3;
                s1_power3_log          <= log_s1_plus_1m2_exp + log_s1_plus_2_exp + "0000000001";
                s3_temp_5              <= s3_temp_4;
                s1_temp_5              <= s1_temp_4;
                s1_s3_flag_3           <= s1_s3_flag_2;
        end if;
end process;
------------------------------------------------------------------------------------------------------------
-- Define processes : (CLK 7)
------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1_pass5  <= "00000001";
                s1_power3_temp   <= "00000001";
                s1_power3_log_1  <= (others => '0');
                s3_temp_6        <= (others => '0');
                s1_temp_6        <= (others => '0');
                s1_s3_flag_4     <= '0';
                hard_input_pass_7<= (others => '0'); 
                soft_input_7     <= (others => (others => '0')); 
        elsif rising_edge(clk) then  
                soft_input_7     <= soft_input_6;
                hard_input_pass_7<= hard_input_pass_6;
                s1_plus_1_pass5  <= s1_plus_1_pass4;
                s1_power3_temp   <= antilog_table(to_integer(unsigned(s1_power3_log)));
                s1_power3_log_1  <= s1_power3_log; -- log(3*s1)
                s3_temp_6        <= s3_temp_5;
                s1_temp_6        <= s1_temp_5;
                s1_s3_flag_4     <= s1_s3_flag_3;
        end if;
end process;
------------------------------------------------------------------------------------------------------------
-- Define processes : (CLK 8)
------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1_pass6  <= "00000001";
                s1_power3        <= "00000001";
                s1_power3_log_2  <= (others => '0');
                s3_temp_7        <= (others => '0');
                s1_temp_7        <= (others => '0');
                s1_power3_exp    <= "000000001";
                s3_temp_6_exp    <= "000000001";
                s1_s3_flag_5     <= '0';
                hard_input_pass_8<= (others => '0'); 
                soft_input_8     <= (others => (others => '0')); 
        elsif rising_edge(clk) then  
                soft_input_8     <= soft_input_7;
                hard_input_pass_8<= hard_input_pass_7;
                s1_plus_1_pass6  <= s1_plus_1_pass5;
                s1_power3        <= s1_power3_temp;
                s1_power3_exp    <= '0' & s1_power3_temp;
                s3_temp_6_exp    <= '0' & s3_temp_6;
                s1_power3_log_2  <= s1_power3_log_1; -- log(3*s1)
                s3_temp_7        <= s3_temp_6;
                s1_temp_7        <= s1_temp_6;
                s1_s3_flag_5     <= s1_s3_flag_4;
        end if;
end process;
------------------------------------------------------------------------------------------------------------
-- Define processes : (CLK 9)
------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1_pass7  <= "00000001";
                s1_power3_1      <= "00000001";
                s1_power3_log_3  <= (others => '0');
                s3_temp_8        <= (others => '0');
                s1_temp_8        <= (others => '0');
                A_index          <= (others => '0');
                s1_s3_flag_6     <= '0';
                s1_power3_s3_flag<= '0';
                hard_input_pass_9<= (others => '0'); 
                soft_input_9     <= (others => (others => '0')); 
        elsif rising_edge(clk) then  
                soft_input_9     <= soft_input_8;
                hard_input_pass_9<= hard_input_pass_8;
                s1_plus_1_pass7  <= s1_plus_1_pass6;
                s1_power3_1      <= s1_power3; -- s1^3
                s1_power3_log_3  <= s1_power3_log_2;
                s3_temp_8        <= s3_temp_7;
                s1_temp_8        <= s1_temp_7;
                A_index          <= s1_power3_exp xor s3_temp_6_exp; -- A calculation
                s1_s3_flag_6     <= s1_s3_flag_5;
                if (s1_power3 = s3_temp_7) then
                        s1_power3_s3_flag <= '1';
                else
                        s1_power3_s3_flag <= '0';
                end if;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 10)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1_pass8    <= "00000001";
                s1_power3_2        <= (others => '0');
                s3_temp_9          <= (others => '0');
                s1_temp_9          <= (others => '0');
                s1_power3_log_4    <= "0000000001";
                log_v              <= (others => '0');
                s1_s3_flag_7       <= '0';
                s1_power3_s3_flag_1<= '0';
                hard_input_pass_10 <= (others => '0'); 
                soft_input_10      <= (others => (others => '0'));
        elsif rising_edge(clk) then  
                soft_input_10      <= soft_input_9;
                hard_input_pass_10 <= hard_input_pass_9;
                s1_plus_1_pass8    <= s1_plus_1_pass7;
                s1_power3_2        <= s1_power3_1;
                s3_temp_9          <= s3_temp_8;
                s1_temp_9          <= s1_temp_8;
                s1_power3_log_4    <= s1_power3_log_3;
                log_v              <= log_table(to_integer(unsigned(A_index)));
                s1_s3_flag_7       <= s1_s3_flag_6;
                s1_power3_s3_flag_1<= s1_power3_s3_flag;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 11)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1_pass9    <= "00000001";
                s1_power3_3        <= (others => '0');
                s3_temp_10         <= (others => '0');
                s1_temp_10         <= (others => '0');
                A_temp             <= 0;
                s1_s3_flag_8       <= '0';
                s1_power3_s3_flag_2<= '0';
                hard_input_pass_11 <= (others => '0'); 
                soft_input_11      <= (others => (others => '0'));
        elsif rising_edge(clk) then  
                soft_input_11      <= soft_input_10;
                hard_input_pass_11 <= hard_input_pass_10;
                s1_plus_1_pass9    <= s1_plus_1_pass8;
                s1_power3_3        <= s1_power3_2;
                s3_temp_10         <= s3_temp_9;
                s1_temp_10         <= s1_temp_9;
                A_temp             <= to_integer(signed(log_v)) - to_integer(unsigned(s1_power3_log_4));
                s1_s3_flag_8       <= s1_s3_flag_7;
                s1_power3_s3_flag_2<= s1_power3_s3_flag_1;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 12)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1_pass10   <= "00000001";
                s1_power3_4        <= (others => '0');
                s3_temp_11         <= (others => '0');
                s1_temp_11         <= (others => '0');
                A                  <= (others => '0');
                s1_s3_flag_9       <= '0';
                s1_power3_s3_flag_3<= '0';
                hard_input_pass_12 <= (others => '0');
                soft_input_12      <= (others => (others => '0')); 
        elsif rising_edge(clk) then 
                soft_input_12      <= soft_input_11; 
                hard_input_pass_12 <= hard_input_pass_11;
                s1_plus_1_pass10   <= s1_plus_1_pass9;
                s1_power3_4        <= s1_power3_3;
                s3_temp_11         <= s3_temp_10;
                s1_temp_11         <= s1_temp_10;
                A                  <= std_logic_vector(to_signed((A_temp + 257),10));
                s1_s3_flag_9       <= s1_s3_flag_8;
                s1_power3_s3_flag_3<= s1_power3_s3_flag_2;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 13)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_plus_1_pass11   <= "00000001";
                s1_power3_5        <= (others => '0');
                s3_temp_12         <= (others => '0');
                s1_temp_12         <= (others => '0');
                xxxc1a             <= (others => '0');
                xxxc2a             <= (others => '0');
                xxxc3a             <= (others => '0');
                s1_s3_flag_10      <= '0';
                s1_power3_s3_flag_4<= '0';
                hard_input_pass_13 <= (others => '0'); 
                soft_input_13      <= (others => (others => '0')); 
        elsif rising_edge(clk) then  
                soft_input_13      <= soft_input_12; 
                hard_input_pass_13 <= hard_input_pass_12;
                s1_plus_1_pass11   <= s1_plus_1_pass10;
                s1_power3_5        <= s1_power3_4;
                s3_temp_12         <= s3_temp_11;
                s1_temp_12         <= s1_temp_11;
                xxxc1a             <= xxxc_1(to_integer(signed(A))); 
                xxxc2a             <= xxxc_2(to_integer(signed(A))); 
                xxxc3a             <= xxxc_3(to_integer(signed(A))); 
                s1_s3_flag_10      <= s1_s3_flag_9;
                s1_power3_s3_flag_4<=s1_power3_s3_flag_3;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 14)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_power3_6        <= (others => '0');
                s3_temp_13         <= (others => '0');
                s1_temp_13         <= (others => '0');
                xxxc2a_1           <= (others => '0');
                xxxc3a_1           <= (others => '0');
                s1_s3_flag_11      <= '0';
                s1_power3_s3_flag_5<= '0';
                log_table_value_s1p<= (others => '0');
                hard_input_pass_14<= (others => '0'); 
                indi_1             <= False;
                indi_2             <= False;
                soft_input_14      <= (others => (others => '0')); 
        elsif rising_edge(clk) then 
                soft_input_14      <= soft_input_13;  
                hard_input_pass_14 <= hard_input_pass_13;
                log_table_value_s1p<= log_table(to_integer(unsigned(s1_plus_1_pass11)));
                s1_power3_6        <= s1_power3_5;
                s3_temp_13         <= s3_temp_12;
                s1_temp_13         <= s1_temp_12;
                xxxc2a_1           <= xxxc2a; 
                xxxc3a_1           <= xxxc3a; 
                s1_s3_flag_11      <= s1_s3_flag_10;
                indi_1             <= (s1_temp_12 /= 0) and (s1_power3_s3_flag_4 = '1');
                indi_2             <= (s1_temp_12 /= 0) and (xxxc1a = 2);
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 15)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                s1_power3_7          <= (others => '0');
                s3_temp_14           <= (others => '0');
                flag_1               <= '0';
                flag_2               <= '0';
                xxxc2a_2             <= (others => '0');
                xxxc3a_2             <= (others => '0');
                s1_s3_flag_12        <= '0';
                s1_power3_s3_flag_6  <= '0';
                log_table_value_s1p_1<= (others => '0');
                hard_input_pass_15   <= (others => '0'); 
                soft_input_15        <= (others => (others => '0')); 
        elsif rising_edge(clk) then 
                soft_input_15        <= soft_input_14;  
                hard_input_pass_15   <= hard_input_pass_14;
                log_table_value_s1p_1<= log_table_value_s1p;
                s1_power3_7          <= s1_power3_6;
                s3_temp_14           <= s3_temp_13;
                xxxc2a_2             <= xxxc2a_1; 
                xxxc3a_2             <= xxxc3a_1; 
                s1_s3_flag_12        <= s1_s3_flag_11;
                if indi_1 then
                        flag_1   <= '1';
                        flag_2   <= '0';
                elsif indi_2 then
                        flag_1   <= '0';
                        flag_2   <= '1';
                else
                        flag_1   <= '0';
                        flag_2   <= '0';
                end if;
        end if;
end process;
------------------------------------------------------------------------------------------------------------
-- Define processes : (CLK 16)
------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                state             <= unable_to_correct_state;
                eh1_temp          <= 255;
                eh2_temp          <= 0;
                eh3_temp          <= 0;
                hard_input_pass_16<= (others => '0'); 
                soft_input_16     <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_16      <= soft_input_15; 
                hard_input_pass_16 <= hard_input_pass_15;
                if s1_s3_flag_12 = '1' then
                        state    <= no_error_state;
                elsif flag_1 = '1' then                                                          -- s1_pass_7 /= 0 and s1_power3_s3_flag_2
                        eh1_temp <= to_integer(unsigned(255 - log_table_value_s1p_1));
                        eh2_temp <= 0;                                                     -- Values for keeping the minus operation functions below
                        eh3_temp <= 0;
                        state    <= one_error_state;
                elsif flag_2 = '1' then                                                           -- s1_pass_7 /= 0 and xxxc1a = 2
                        eh1_temp <= 255;
                        eh2_temp <= to_integer(unsigned(xxxc2a_2 + log_table_value_s1p_1)); -- xxxc(A,2)+log_table(S1+1)
                        eh3_temp <= to_integer(unsigned(xxxc3a_2 + log_table_value_s1p_1));
                        state    <= two_error_state;
                else
                        eh1_temp <= 255;                                                    -- When nothing happens, this is the default value
                        eh2_temp <= 0;
                        eh3_temp <= 0;
                        state    <= unable_to_correct_state;
                end if;
        end if;
end process;
----------------------------------------------------------------------------------------------------------------
------ Define processes : (CLK 17)
----------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                next_state        <= unable_to_correct_state;
                eh1_n1            <= 255;
                eh1_n2            <= 255;
                hard_input_f      <= (others => '0');
                eh1               <= 256;
                eh2               <= 256;
                eh3               <= 256;
                soft_input_17     <= (others => (others => '0'));
        elsif rising_edge(clk) then  
                soft_input_17     <= soft_input_16;
                next_state        <= state;
                hard_input_f      <= hard_input_pass_16;
                eh1_n1            <= eh1_temp - 1;                   -- eh1 - 1        
                eh1_n2            <= eh1_temp - 2;                   -- eh1 - 2    
                eh1               <= eh1_temp;                       -- eh1
                if eh2_temp > 509 then                               -- Need to bring this value back to range, eh2 and eh3 are ready, all in integer
                        eh2 <= 765 - eh2_temp;
                elsif eh2_temp > 254 then                            -- 
                        eh2 <= 510 - eh2_temp;
                else
                        eh2 <= 255 - eh2_temp;    
                end if;
                if eh3_temp > 509 then
                        eh3 <= 765 - eh3_temp;
                elsif eh3_temp > 254 then
                        eh3 <= 510 - eh3_temp;
                else
                        eh3 <= 255 - eh3_temp;    
                end if;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 18)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_temp  <= (others => '0');
                eh1_pass          <= 255;
                eh2_pass          <= 255;
                eh3_pass          <= 255;
                eh1_pass_n1       <= 255;
                eh1_pass_n2       <= 255;
                eh2_pass_n1       <= 255;
                eh3_pass_n1       <= 255; 
                next_state_1      <= unable_to_correct_state;  
                soft_input_18     <= (others => (others => '0'));        
        elsif rising_edge(clk) then 
                soft_input_18     <= soft_input_17;
                next_state_1      <= next_state;
                eh1_pass_n1       <= eh1_n1;
                eh1_pass_n2       <= eh1_n2;
                eh1_pass          <= eh1;
                eh2_pass          <= eh2;
                eh2_pass_n1       <= eh2 - 1;
                eh3_pass          <= eh3;
                eh3_pass_n1       <= eh3 - 1;      -- prepare for next clock cycle
                hard_output_temp  <= hard_input_f; -- keep on passing the hard input
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 19)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                next_state_2             <= unable_to_correct_state;  
                hard_output_error_1      <= '0';
                hard_output_error_2      <= '0';
                hard_output_error_3      <= '0';
                hard_output_error_rest_1 <= (others => '0');
                eh1_pass_1               <= 255;
                eh2_pass_1               <= 255;
                eh3_pass_1               <= 255;
                eh1_pass_n1_1            <= 255;
                eh2_pass_n1_1            <= 255;
                eh3_pass_n1_1            <= 255;
                soft_input_19            <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_19            <= soft_input_18;
                next_state_2             <= next_state_1;  
                hard_output_error_1      <= not hard_output_temp(eh1_pass_n1);
                hard_output_error_2      <= not hard_output_temp(eh2_pass_n1);
                hard_output_error_3      <= not hard_output_temp(eh3_pass_n1);
                hard_output_error_rest_1 <= hard_output_temp; -- original input
                eh1_pass_1               <= eh1_pass;
                eh2_pass_1               <= eh2_pass;
                eh3_pass_1               <= eh3_pass;
                eh1_pass_n1_1            <= eh1_pass_n1;
                eh2_pass_n1_1            <= eh2_pass_n1;
                eh3_pass_n1_1            <= eh3_pass_n1;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 20)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                error_position_temp(0)          <= -1;
                error_position_temp(1)          <= -1;
                error_position_temp(2)          <= -1;
                hard_output_error_rest_2        <= (others => '0');
                corrections_temp                <= "000";
                soft_input_20                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_20                   <= soft_input_19;
                case next_state_2 is
                        when no_error_state =>
                                corrections_temp                        <= "000";
                                hard_output_error_rest_2                <= hard_output_error_rest_1; -- Unable to correct, input goes to output 
                                error_position_temp(0)                  <= -1;
                                error_position_temp(1)                  <= -1;
                                error_position_temp(2)                  <= -1;
                        when one_error_state =>
                                corrections_temp                        <= "001";
                                hard_output_error_rest_2                <= hard_output_error_rest_1;
                                hard_output_error_rest_2(eh1_pass_n1_1) <= hard_output_error_1;
                                error_position_temp(0)                  <= eh1_pass_1;
                                error_position_temp(1)                  <= -1;
                                error_position_temp(2)                  <= -1;
                        when two_error_state =>
                                corrections_temp                        <= "010";
                                hard_output_error_rest_2                <= hard_output_error_rest_1;
                                hard_output_error_rest_2(eh2_pass_n1_1) <= hard_output_error_2;
                                hard_output_error_rest_2(eh3_pass_n1_1) <= hard_output_error_3;
                                error_position_temp(0)                  <= eh2_pass_1;
                                error_position_temp(1)                  <= eh3_pass_1;
                                error_position_temp(2)                  <= -1;                       -- reserved for parity error
                        when unable_to_correct_state =>
                                corrections_temp                        <= "100";
                                hard_output_error_rest_2                <= hard_output_error_rest_1; -- Unable to correct, input goes to output   
                                error_position_temp(0)                  <= -1;
                                error_position_temp(1)                  <= -1;
                                error_position_temp(2)                  <= -1;      
                end case; 
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 21) Start calculating sum
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_3        <= (others => '0');
                error_position_temp_1(0)        <= -1;
                error_position_temp_1(1)        <= -1;
                error_position_temp_1(2)        <= -1;
                corrections_temp_1              <= "000";
                sum_1_1                         <= (others => '0');
                sum_1_2                         <= (others => '0');
                sum_1_3                         <= (others => '0');
                sum_1_4                         <= (others => '0');
                soft_input_21                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                --------------------------------------------------------------------------------------------------------------
                -- Output can be tested here
                --corrections    <= corrections_temp;
                --error_position <= error_position_temp;
                --hard_output    <= hard_output_error_rest_2;
                --sum            <= sum_16_temp_3;
                --------------------------------------------------------------------------------------------------------------
                soft_input_21                   <= soft_input_20;
                hard_output_error_rest_3        <= hard_output_error_rest_2;                            -- pass the corrected data
                error_position_temp_1           <= error_position_temp;                                 -- passing the error position
                corrections_temp_1              <= corrections_temp;                                    -- passing the correction number
                sum_1_1                         <= ("00000000"&hard_output_error_rest_2(0)) + ("00000000"&hard_output_error_rest_2(1)) + ("00000000"&hard_output_error_rest_2(2)) + ("00000000"&hard_output_error_rest_2(3));
                sum_1_2                         <= ("00000000"&hard_output_error_rest_2(4)) + ("00000000"&hard_output_error_rest_2(5)) + ("00000000"&hard_output_error_rest_2(6)) + ("00000000"&hard_output_error_rest_2(7));
                sum_1_3                         <= ("00000000"&hard_output_error_rest_2(8)) + ("00000000"&hard_output_error_rest_2(9)) + ("00000000"&hard_output_error_rest_2(10)) + ("00000000"&hard_output_error_rest_2(11));
                sum_1_4                         <= ("00000000"&hard_output_error_rest_2(12)) + ("00000000"&hard_output_error_rest_2(13)) + ("00000000"&hard_output_error_rest_2(14)) + ("00000000"&hard_output_error_rest_2(15));
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 22)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_4        <= (others => '0');
                error_position_temp_2(0)        <= -1;
                error_position_temp_2(1)        <= -1;
                error_position_temp_2(2)        <= -1;
                corrections_temp_2              <= "000";
                sum_2_1                         <= (others => '0');
                sum_2_2                         <= (others => '0');
                sum_2_3                         <= (others => '0');
                sum_2_4                         <= (others => '0');
                sum_2_5                         <= (others => '0');
                soft_input_22                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_22                   <= soft_input_21;
                hard_output_error_rest_4        <= hard_output_error_rest_3;                            -- pass the corrected data
                error_position_temp_2           <= error_position_temp_1;                                 -- passing the error position
                corrections_temp_2              <= corrections_temp_1;                                    -- passing the correction number
                sum_2_1                         <= ("00000000"&hard_output_error_rest_3(16)) + ("00000000"&hard_output_error_rest_3(17)) + ("00000000"&hard_output_error_rest_3(18)) + ("00000000"&hard_output_error_rest_3(19));
                sum_2_2                         <= ("00000000"&hard_output_error_rest_3(20)) + ("00000000"&hard_output_error_rest_3(21)) + ("00000000"&hard_output_error_rest_3(22)) + ("00000000"&hard_output_error_rest_3(23));
                sum_2_3                         <= ("00000000"&hard_output_error_rest_3(24)) + ("00000000"&hard_output_error_rest_3(25)) + ("00000000"&hard_output_error_rest_3(26)) + ("00000000"&hard_output_error_rest_3(27));
                sum_2_4                         <= ("00000000"&hard_output_error_rest_3(28)) + ("00000000"&hard_output_error_rest_3(29)) + ("00000000"&hard_output_error_rest_3(30)) + ("00000000"&hard_output_error_rest_3(31));
                sum_2_5                         <= sum_1_1 + sum_1_2 + sum_1_3 + sum_1_4;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 23)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_5        <= (others => '0');
                error_position_temp_3(0)        <= -1;
                error_position_temp_3(1)        <= -1;
                error_position_temp_3(2)        <= -1;
                corrections_temp_3              <= "000";
                sum_3_1                         <= (others => '0');
                sum_3_2                         <= (others => '0');
                sum_3_3                         <= (others => '0');
                sum_3_4                         <= (others => '0');
                sum_3_5                         <= (others => '0');
                soft_input_23                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_23                   <= soft_input_22;
                hard_output_error_rest_5        <= hard_output_error_rest_4;                              -- pass the corrected data
                error_position_temp_3           <= error_position_temp_2;                                 -- passing the error position
                corrections_temp_3              <= corrections_temp_2;                                    -- passing the correction number
                sum_3_1                         <= ("00000000"&hard_output_error_rest_4(32)) + ("00000000"&hard_output_error_rest_4(33)) + ("00000000"&hard_output_error_rest_4(34)) + ("00000000"&hard_output_error_rest_4(35));
                sum_3_2                         <= ("00000000"&hard_output_error_rest_4(36)) + ("00000000"&hard_output_error_rest_4(37)) + ("00000000"&hard_output_error_rest_4(38)) + ("00000000"&hard_output_error_rest_4(39));
                sum_3_3                         <= ("00000000"&hard_output_error_rest_4(40)) + ("00000000"&hard_output_error_rest_4(41)) + ("00000000"&hard_output_error_rest_4(42)) + ("00000000"&hard_output_error_rest_4(43));
                sum_3_4                         <= ("00000000"&hard_output_error_rest_4(44)) + ("00000000"&hard_output_error_rest_4(45)) + ("00000000"&hard_output_error_rest_4(46)) + ("00000000"&hard_output_error_rest_4(47));
                sum_3_5                         <= sum_2_1 + sum_2_2 + sum_2_3 + sum_2_4 + sum_2_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 24)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_6        <= (others => '0');
                error_position_temp_4(0)        <= -1;
                error_position_temp_4(1)        <= -1;
                error_position_temp_4(2)        <= -1;
                corrections_temp_4              <= "000";
                sum_4_1                         <= (others => '0');
                sum_4_2                         <= (others => '0');
                sum_4_3                         <= (others => '0');
                sum_4_4                         <= (others => '0');
                sum_4_5                         <= (others => '0');
                soft_input_24                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_24                   <= soft_input_23;
                hard_output_error_rest_6        <= hard_output_error_rest_5;                              -- pass the corrected data
                error_position_temp_4           <= error_position_temp_3;                                 -- passing the error position
                corrections_temp_4              <= corrections_temp_3;                                    -- passing the correction number
                sum_4_1                         <= ("00000000"&hard_output_error_rest_5(48)) + ("00000000"&hard_output_error_rest_5(49)) + ("00000000"&hard_output_error_rest_5(50)) + ("00000000"&hard_output_error_rest_5(51));
                sum_4_2                         <= ("00000000"&hard_output_error_rest_5(52)) + ("00000000"&hard_output_error_rest_5(53)) + ("00000000"&hard_output_error_rest_5(54)) + ("00000000"&hard_output_error_rest_5(55));
                sum_4_3                         <= ("00000000"&hard_output_error_rest_5(56)) + ("00000000"&hard_output_error_rest_5(57)) + ("00000000"&hard_output_error_rest_5(58)) + ("00000000"&hard_output_error_rest_5(59));
                sum_4_4                         <= ("00000000"&hard_output_error_rest_5(60)) + ("00000000"&hard_output_error_rest_5(61)) + ("00000000"&hard_output_error_rest_5(62)) + ("00000000"&hard_output_error_rest_5(63));
                sum_4_5                         <= sum_3_1 + sum_3_2 + sum_3_3 + sum_3_4 + sum_3_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 25)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_7        <= (others => '0');
                error_position_temp_5(0)        <= -1;
                error_position_temp_5(1)        <= -1;
                error_position_temp_5(2)        <= -1;
                corrections_temp_5              <= "000";
                sum_5_1                         <= (others => '0');
                sum_5_2                         <= (others => '0');
                sum_5_3                         <= (others => '0');
                sum_5_4                         <= (others => '0');
                sum_5_5                         <= (others => '0');
                soft_input_25                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_25                   <= soft_input_24;
                hard_output_error_rest_7        <= hard_output_error_rest_6;                              -- pass the corrected data
                error_position_temp_5           <= error_position_temp_4;                                 -- passing the error position
                corrections_temp_5              <= corrections_temp_4;                                    -- passing the correction number
                sum_5_1                         <= ("00000000"&hard_output_error_rest_6(64)) + ("00000000"&hard_output_error_rest_6(65)) + ("00000000"&hard_output_error_rest_6(66)) + ("00000000"&hard_output_error_rest_6(67));
                sum_5_2                         <= ("00000000"&hard_output_error_rest_6(68)) + ("00000000"&hard_output_error_rest_6(69)) + ("00000000"&hard_output_error_rest_6(70)) + ("00000000"&hard_output_error_rest_6(71));
                sum_5_3                         <= ("00000000"&hard_output_error_rest_6(72)) + ("00000000"&hard_output_error_rest_6(73)) + ("00000000"&hard_output_error_rest_6(74)) + ("00000000"&hard_output_error_rest_6(75));
                sum_5_4                         <= ("00000000"&hard_output_error_rest_6(76)) + ("00000000"&hard_output_error_rest_6(77)) + ("00000000"&hard_output_error_rest_6(78)) + ("00000000"&hard_output_error_rest_6(79));
                sum_5_5                         <= sum_4_1 + sum_4_2 + sum_4_3 + sum_4_4 + sum_4_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 26)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_8        <= (others => '0');
                error_position_temp_6(0)        <= -1;
                error_position_temp_6(1)        <= -1;
                error_position_temp_6(2)        <= -1;
                corrections_temp_6              <= "000";
                sum_6_1                         <= (others => '0');
                sum_6_2                         <= (others => '0');
                sum_6_3                         <= (others => '0');
                sum_6_4                         <= (others => '0');
                sum_6_5                         <= (others => '0');
                soft_input_26                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_26                   <= soft_input_25;
                hard_output_error_rest_8        <= hard_output_error_rest_7;                              -- pass the corrected data
                error_position_temp_6           <= error_position_temp_5;                                 -- passing the error position
                corrections_temp_6              <= corrections_temp_5;                                    -- passing the correction number
                sum_6_1                         <= ("00000000"&hard_output_error_rest_7(80)) + ("00000000"&hard_output_error_rest_7(81)) + ("00000000"&hard_output_error_rest_7(82)) + ("00000000"&hard_output_error_rest_7(83));
                sum_6_2                         <= ("00000000"&hard_output_error_rest_7(84)) + ("00000000"&hard_output_error_rest_7(85)) + ("00000000"&hard_output_error_rest_7(86)) + ("00000000"&hard_output_error_rest_7(87));
                sum_6_3                         <= ("00000000"&hard_output_error_rest_7(88)) + ("00000000"&hard_output_error_rest_7(89)) + ("00000000"&hard_output_error_rest_7(90)) + ("00000000"&hard_output_error_rest_7(91));
                sum_6_4                         <= ("00000000"&hard_output_error_rest_7(92)) + ("00000000"&hard_output_error_rest_7(93)) + ("00000000"&hard_output_error_rest_7(94)) + ("00000000"&hard_output_error_rest_7(95));
                sum_6_5                         <= sum_5_1 + sum_5_2 + sum_5_3 + sum_5_4 + sum_5_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 27)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_9        <= (others => '0');
                error_position_temp_7(0)        <= -1;
                error_position_temp_7(1)        <= -1;
                error_position_temp_7(2)        <= -1;
                corrections_temp_7              <= "000";
                sum_7_1                         <= (others => '0');
                sum_7_2                         <= (others => '0');
                sum_7_3                         <= (others => '0');
                sum_7_4                         <= (others => '0');
                sum_7_5                         <= (others => '0');
                soft_input_27                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_27                   <= soft_input_26;
                hard_output_error_rest_9        <= hard_output_error_rest_8;                              -- pass the corrected data
                error_position_temp_7           <= error_position_temp_6;                                 -- passing the error position
                corrections_temp_7              <= corrections_temp_6;                                    -- passing the correction number
                sum_7_1                         <= ("00000000"&hard_output_error_rest_8(96)) + ("00000000"&hard_output_error_rest_8(97)) + ("00000000"&hard_output_error_rest_8(98)) + ("00000000"&hard_output_error_rest_8(99));
                sum_7_2                         <= ("00000000"&hard_output_error_rest_8(100)) + ("00000000"&hard_output_error_rest_8(101)) + ("00000000"&hard_output_error_rest_8(102)) + ("00000000"&hard_output_error_rest_8(103));
                sum_7_3                         <= ("00000000"&hard_output_error_rest_8(104)) + ("00000000"&hard_output_error_rest_8(105)) + ("00000000"&hard_output_error_rest_8(106)) + ("00000000"&hard_output_error_rest_8(107));
                sum_7_4                         <= ("00000000"&hard_output_error_rest_8(108)) + ("00000000"&hard_output_error_rest_8(109)) + ("00000000"&hard_output_error_rest_8(110)) + ("00000000"&hard_output_error_rest_8(111));
                sum_7_5                         <= sum_6_1 + sum_6_2 + sum_6_3 + sum_6_4 + sum_6_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 28)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_10       <= (others => '0');
                error_position_temp_8(0)        <= -1;
                error_position_temp_8(1)        <= -1;
                error_position_temp_8(2)        <= -1;
                corrections_temp_8              <= "000";
                sum_8_1                         <= (others => '0');
                sum_8_2                         <= (others => '0');
                sum_8_3                         <= (others => '0');
                sum_8_4                         <= (others => '0');
                sum_8_5                         <= (others => '0');
                soft_input_28                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_28                   <= soft_input_27;
                hard_output_error_rest_10       <= hard_output_error_rest_9;                              -- pass the corrected data
                error_position_temp_8           <= error_position_temp_7;                                 -- passing the error position
                corrections_temp_8              <= corrections_temp_7;                                    -- passing the correction number
                sum_8_1                         <= ("00000000"&hard_output_error_rest_9(112)) + ("00000000"&hard_output_error_rest_9(113)) + ("00000000"&hard_output_error_rest_9(114)) + ("00000000"&hard_output_error_rest_9(115));
                sum_8_2                         <= ("00000000"&hard_output_error_rest_9(116)) + ("00000000"&hard_output_error_rest_9(117)) + ("00000000"&hard_output_error_rest_9(118)) + ("00000000"&hard_output_error_rest_9(119));
                sum_8_3                         <= ("00000000"&hard_output_error_rest_9(120)) + ("00000000"&hard_output_error_rest_9(121)) + ("00000000"&hard_output_error_rest_9(122)) + ("00000000"&hard_output_error_rest_9(123));
                sum_8_4                         <= ("00000000"&hard_output_error_rest_9(124)) + ("00000000"&hard_output_error_rest_9(125)) + ("00000000"&hard_output_error_rest_9(126)) + ("00000000"&hard_output_error_rest_9(127));
                sum_8_5                         <= sum_7_1 + sum_7_2 + sum_7_3 + sum_7_4 + sum_7_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 29)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_11       <= (others => '0');
                error_position_temp_9(0)        <= -1;
                error_position_temp_9(1)        <= -1;
                error_position_temp_9(2)        <= -1;
                corrections_temp_9              <= "000";
                sum_9_1                         <= (others => '0');
                sum_9_2                         <= (others => '0');
                sum_9_3                         <= (others => '0');
                sum_9_4                         <= (others => '0');
                sum_9_5                         <= (others => '0');
                soft_input_29                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_29                   <= soft_input_28;
                hard_output_error_rest_11       <= hard_output_error_rest_10;                             -- pass the corrected data
                error_position_temp_9           <= error_position_temp_8;                                 -- passing the error position
                corrections_temp_9              <= corrections_temp_8;                                    -- passing the correction number
                sum_9_1                         <= ("00000000"&hard_output_error_rest_10(128)) + ("00000000"&hard_output_error_rest_10(129)) + ("00000000"&hard_output_error_rest_10(130)) + ("00000000"&hard_output_error_rest_10(131));
                sum_9_2                         <= ("00000000"&hard_output_error_rest_10(132)) + ("00000000"&hard_output_error_rest_10(133)) + ("00000000"&hard_output_error_rest_10(134)) + ("00000000"&hard_output_error_rest_10(135));
                sum_9_3                         <= ("00000000"&hard_output_error_rest_10(136)) + ("00000000"&hard_output_error_rest_10(137)) + ("00000000"&hard_output_error_rest_10(138)) + ("00000000"&hard_output_error_rest_10(139));
                sum_9_4                         <= ("00000000"&hard_output_error_rest_10(140)) + ("00000000"&hard_output_error_rest_10(141)) + ("00000000"&hard_output_error_rest_10(142)) + ("00000000"&hard_output_error_rest_10(143));
                sum_9_5                         <= sum_8_1 + sum_8_2 + sum_8_3 + sum_8_4 + sum_8_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 30)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_12        <= (others => '0');
                error_position_temp_10(0)        <= -1;
                error_position_temp_10(1)        <= -1;
                error_position_temp_10(2)        <= -1;
                corrections_temp_10              <= "000";
                sum_10_1                         <= (others => '0');
                sum_10_2                         <= (others => '0');
                sum_10_3                         <= (others => '0');
                sum_10_4                         <= (others => '0');
                sum_10_5                         <= (others => '0');
                soft_input_30                    <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_30                    <= soft_input_29;
                hard_output_error_rest_12        <= hard_output_error_rest_11;                             -- pass the corrected data
                error_position_temp_10           <= error_position_temp_9;                                 -- passing the error position
                corrections_temp_10              <= corrections_temp_9;                                    -- passing the correction number
                sum_10_1                         <= ("00000000"&hard_output_error_rest_11(144)) + ("00000000"&hard_output_error_rest_11(145)) + ("00000000"&hard_output_error_rest_11(146)) + ("00000000"&hard_output_error_rest_11(147));
                sum_10_2                         <= ("00000000"&hard_output_error_rest_11(148)) + ("00000000"&hard_output_error_rest_11(149)) + ("00000000"&hard_output_error_rest_11(150)) + ("00000000"&hard_output_error_rest_11(151));
                sum_10_3                         <= ("00000000"&hard_output_error_rest_11(152)) + ("00000000"&hard_output_error_rest_11(153)) + ("00000000"&hard_output_error_rest_11(154)) + ("00000000"&hard_output_error_rest_11(155));
                sum_10_4                         <= ("00000000"&hard_output_error_rest_11(156)) + ("00000000"&hard_output_error_rest_11(157)) + ("00000000"&hard_output_error_rest_11(158)) + ("00000000"&hard_output_error_rest_11(159));
                sum_10_5                         <= sum_9_1 + sum_9_2 + sum_9_3 + sum_9_4 + sum_9_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 31)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_13        <= (others => '0');
                error_position_temp_11(0)        <= -1;
                error_position_temp_11(1)        <= -1;
                error_position_temp_11(2)        <= -1;
                corrections_temp_11              <= "000";
                sum_11_1                         <= (others => '0');
                sum_11_2                         <= (others => '0');
                sum_11_3                         <= (others => '0');
                sum_11_4                         <= (others => '0');
                sum_11_5                         <= (others => '0');
                soft_input_31                    <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_31                    <= soft_input_30;
                hard_output_error_rest_13        <= hard_output_error_rest_12;                              -- pass the corrected data
                error_position_temp_11           <= error_position_temp_10;                                 -- passing the error position
                corrections_temp_11              <= corrections_temp_10;                                    -- passing the correction number
                sum_11_1                         <= ("00000000"&hard_output_error_rest_12(160)) + ("00000000"&hard_output_error_rest_12(161)) + ("00000000"&hard_output_error_rest_12(162)) + ("00000000"&hard_output_error_rest_12(163));
                sum_11_2                         <= ("00000000"&hard_output_error_rest_12(164)) + ("00000000"&hard_output_error_rest_12(165)) + ("00000000"&hard_output_error_rest_12(166)) + ("00000000"&hard_output_error_rest_12(167));
                sum_11_3                         <= ("00000000"&hard_output_error_rest_12(168)) + ("00000000"&hard_output_error_rest_12(169)) + ("00000000"&hard_output_error_rest_12(170)) + ("00000000"&hard_output_error_rest_12(171));
                sum_11_4                         <= ("00000000"&hard_output_error_rest_12(172)) + ("00000000"&hard_output_error_rest_12(173)) + ("00000000"&hard_output_error_rest_12(174)) + ("00000000"&hard_output_error_rest_12(175));
                sum_11_5                         <= sum_10_1 + sum_10_2 + sum_10_3 + sum_10_4 + sum_10_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 32)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_14        <= (others => '0');
                error_position_temp_12(0)        <= -1;
                error_position_temp_12(1)        <= -1;
                error_position_temp_12(2)        <= -1;
                corrections_temp_12              <= "000";
                sum_12_1                         <= (others => '0');
                sum_12_2                         <= (others => '0');
                sum_12_3                         <= (others => '0');
                sum_12_4                         <= (others => '0');
                sum_12_5                         <= (others => '0');
                soft_input_32                    <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_32                    <= soft_input_31;
                hard_output_error_rest_14        <= hard_output_error_rest_13;                              -- pass the corrected data
                error_position_temp_12           <= error_position_temp_11;                                 -- passing the error position
                corrections_temp_12              <= corrections_temp_11;                                    -- passing the correction number
                sum_12_1                         <= ("00000000"&hard_output_error_rest_13(176)) + ("00000000"&hard_output_error_rest_13(177)) + ("00000000"&hard_output_error_rest_13(178)) + ("00000000"&hard_output_error_rest_13(179));
                sum_12_2                         <= ("00000000"&hard_output_error_rest_13(180)) + ("00000000"&hard_output_error_rest_13(181)) + ("00000000"&hard_output_error_rest_13(182)) + ("00000000"&hard_output_error_rest_13(183));
                sum_12_3                         <= ("00000000"&hard_output_error_rest_13(184)) + ("00000000"&hard_output_error_rest_13(185)) + ("00000000"&hard_output_error_rest_13(186)) + ("00000000"&hard_output_error_rest_13(187));
                sum_12_4                         <= ("00000000"&hard_output_error_rest_13(188)) + ("00000000"&hard_output_error_rest_13(189)) + ("00000000"&hard_output_error_rest_13(190)) + ("00000000"&hard_output_error_rest_13(191));
                sum_12_5                         <= sum_11_1 + sum_11_2 + sum_11_3 + sum_11_4 + sum_11_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 33)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_15        <= (others => '0');
                error_position_temp_13(0)        <= -1;
                error_position_temp_13(1)        <= -1;
                error_position_temp_13(2)        <= -1;
                corrections_temp_13              <= "000";
                sum_13_1                         <= (others => '0');
                sum_13_2                         <= (others => '0');
                sum_13_3                         <= (others => '0');
                sum_13_4                         <= (others => '0');
                sum_13_5                         <= (others => '0');
                soft_input_33                    <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_33                    <= soft_input_32;
                hard_output_error_rest_15        <= hard_output_error_rest_14;                              -- pass the corrected data
                error_position_temp_13           <= error_position_temp_12;                                 -- passing the error position
                corrections_temp_13              <= corrections_temp_12;                                    -- passing the correction number
                sum_13_1                         <= ("00000000"&hard_output_error_rest_14(192)) + ("00000000"&hard_output_error_rest_14(193)) + ("00000000"&hard_output_error_rest_14(194)) + ("00000000"&hard_output_error_rest_14(195));
                sum_13_2                         <= ("00000000"&hard_output_error_rest_14(196)) + ("00000000"&hard_output_error_rest_14(197)) + ("00000000"&hard_output_error_rest_14(198)) + ("00000000"&hard_output_error_rest_14(199));
                sum_13_3                         <= ("00000000"&hard_output_error_rest_14(200)) + ("00000000"&hard_output_error_rest_14(201)) + ("00000000"&hard_output_error_rest_14(202)) + ("00000000"&hard_output_error_rest_14(203));
                sum_13_4                         <= ("00000000"&hard_output_error_rest_14(204)) + ("00000000"&hard_output_error_rest_14(205)) + ("00000000"&hard_output_error_rest_14(206)) + ("00000000"&hard_output_error_rest_14(207));
                sum_13_5                         <= sum_12_1 + sum_12_2 + sum_12_3 + sum_12_4 + sum_12_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 34)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_16        <= (others => '0');
                error_position_temp_14(0)        <= -1;
                error_position_temp_14(1)        <= -1;
                error_position_temp_14(2)        <= -1;
                corrections_temp_14              <= "000";
                sum_14_1                         <= (others => '0');
                sum_14_2                         <= (others => '0');
                sum_14_3                         <= (others => '0');
                sum_14_4                         <= (others => '0');
                sum_14_5                         <= (others => '0');
                soft_input_34                    <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_34                    <= soft_input_33;
                hard_output_error_rest_16        <= hard_output_error_rest_15;                              -- pass the corrected data
                error_position_temp_14           <= error_position_temp_13;                                 -- passing the error position
                corrections_temp_14              <= corrections_temp_13;                                    -- passing the correction number
                sum_14_1                         <= ("00000000"&hard_output_error_rest_15(208)) + ("00000000"&hard_output_error_rest_15(209)) + ("00000000"&hard_output_error_rest_15(210)) + ("00000000"&hard_output_error_rest_15(211));
                sum_14_2                         <= ("00000000"&hard_output_error_rest_15(212)) + ("00000000"&hard_output_error_rest_15(213)) + ("00000000"&hard_output_error_rest_15(214)) + ("00000000"&hard_output_error_rest_15(215));
                sum_14_3                         <= ("00000000"&hard_output_error_rest_15(216)) + ("00000000"&hard_output_error_rest_15(217)) + ("00000000"&hard_output_error_rest_15(218)) + ("00000000"&hard_output_error_rest_15(219));
                sum_14_4                         <= ("00000000"&hard_output_error_rest_15(220)) + ("00000000"&hard_output_error_rest_15(221)) + ("00000000"&hard_output_error_rest_15(222)) + ("00000000"&hard_output_error_rest_15(223));
                sum_14_5                         <= sum_13_1 + sum_13_2 + sum_13_3 + sum_13_4 + sum_13_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 35)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_17        <= (others => '0');
                error_position_temp_15(0)        <= -1;
                error_position_temp_15(1)        <= -1;
                error_position_temp_15(2)        <= -1;
                corrections_temp_15              <= "000";
                sum_15_1                         <= (others => '0');
                sum_15_2                         <= (others => '0');
                sum_15_3                         <= (others => '0');
                sum_15_4                         <= (others => '0');
                sum_15_5                         <= (others => '0');
                soft_input_35                    <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_35                    <= soft_input_34;
                hard_output_error_rest_17        <= hard_output_error_rest_16;                              -- pass the corrected data
                error_position_temp_15           <= error_position_temp_14;                                 -- passing the error position
                corrections_temp_15              <= corrections_temp_14;                                    -- passing the correction number
                sum_15_1                         <= ("00000000"&hard_output_error_rest_16(224)) + ("00000000"&hard_output_error_rest_16(225)) + ("00000000"&hard_output_error_rest_16(226)) + ("00000000"&hard_output_error_rest_16(227));
                sum_15_2                         <= ("00000000"&hard_output_error_rest_16(228)) + ("00000000"&hard_output_error_rest_16(229)) + ("00000000"&hard_output_error_rest_16(230)) + ("00000000"&hard_output_error_rest_16(231));
                sum_15_3                         <= ("00000000"&hard_output_error_rest_16(232)) + ("00000000"&hard_output_error_rest_16(233)) + ("00000000"&hard_output_error_rest_16(234)) + ("00000000"&hard_output_error_rest_16(235));
                sum_15_4                         <= ("00000000"&hard_output_error_rest_16(236)) + ("00000000"&hard_output_error_rest_16(237)) + ("00000000"&hard_output_error_rest_16(238)) + ("00000000"&hard_output_error_rest_16(239));
                sum_15_5                         <= sum_14_1 + sum_14_2 + sum_14_3 + sum_14_4 + sum_14_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 36)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_18        <= (others => '0');
                error_position_temp_16(0)        <= -1;
                error_position_temp_16(1)        <= -1;
                error_position_temp_16(2)        <= -1;
                corrections_temp_16              <= "000";
                sum_16_1                         <= (others => '0');
                sum_16_2                         <= (others => '0');
                sum_16_3                         <= (others => '0');
                sum_16_4                         <= (others => '0');
                sum_16_5                         <= (others => '0');
                soft_input_36                    <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_36                    <= soft_input_35;
                hard_output_error_rest_18        <= hard_output_error_rest_17;                              -- pass the corrected data
                error_position_temp_16           <= error_position_temp_15;                                 -- passing the error position
                corrections_temp_16              <= corrections_temp_15;                                    -- passing the correction number
                sum_16_1                         <= ("00000000"&hard_output_error_rest_17(240)) + ("00000000"&hard_output_error_rest_17(241)) + ("00000000"&hard_output_error_rest_17(242)) + ("00000000"&hard_output_error_rest_17(243));
                sum_16_2                         <= ("00000000"&hard_output_error_rest_17(244)) + ("00000000"&hard_output_error_rest_17(245)) + ("00000000"&hard_output_error_rest_17(246)) + ("00000000"&hard_output_error_rest_17(247));
                sum_16_3                         <= ("00000000"&hard_output_error_rest_17(248)) + ("00000000"&hard_output_error_rest_17(249)) + ("00000000"&hard_output_error_rest_17(250)) + ("00000000"&hard_output_error_rest_17(251));
                sum_16_4                         <= ("00000000"&hard_output_error_rest_17(252)) + ("00000000"&hard_output_error_rest_17(253)) + ("00000000"&hard_output_error_rest_17(254));
                sum_16_5                         <= sum_15_1 + sum_15_2 + sum_15_3 + sum_15_4 + sum_15_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 36)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_19        <= (others => '0');
                error_position_temp_17(0)        <= -1;
                error_position_temp_17(1)        <= -1;
                error_position_temp_17(2)        <= -1;
                corrections_temp_17              <= "000";
                sum_16_temp_1                    <= (others => '0');
                soft_input_37                    <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_37                    <= soft_input_36;
                hard_output_error_rest_19        <= hard_output_error_rest_18;                              -- pass the corrected data
                error_position_temp_17           <= error_position_temp_16;                                 -- passing the error position
                corrections_temp_17              <= corrections_temp_16;                                    -- passing the correction number
                sum_16_temp_1                    <= sum_16_1 + sum_16_2 + sum_16_3 + sum_16_4 + sum_16_5;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 21) Start checking the last bit
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                indi_3                          <= False;
                hard_output_error_rest_20       <= (others => '0');
                last_bit                        <= '0';
                error_position_temp_18(0)       <= -1;
                error_position_temp_18(1)       <= -1;
                error_position_temp_18(2)       <= -1;
                corrections_temp_18             <= "000";
                soft_input_38                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                --------------------------------------------------------------------------------------------------------------
                -- Output can be tested here
                --corrections    <= corrections_temp;
                --error_position <= error_position_temp;
                --hard_output    <= hard_output_error_rest_2;
                --sum            <= sum_16_temp_3;
                --------------------------------------------------------------------------------------------------------------
                soft_input_38                   <= soft_input_37;
                indi_3                          <= (hard_output_error_rest_19(255) /= sum_16_temp_1(0)); -- (Decoded(256) ~= mod(sum(Decoded(1:255)),2)) 
                hard_output_error_rest_20       <= hard_output_error_rest_19;                            -- pass the corrected data
                last_bit                        <= not hard_output_error_rest_19(255);                   -- flip it anyway, store it here
                error_position_temp_18          <= error_position_temp_17;                               -- passing the error position
                corrections_temp_18             <= corrections_temp_17;                                  -- passing the correction number
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 22)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                indi_4                          <= False;
                hard_output_error_rest_21       <= (others => '0');
                last_bit_1                      <= '0';
                error_position_temp_19(0)       <= -1;
                error_position_temp_19(1)       <= -1;
                error_position_temp_19(2)       <= -1;
                corrections_temp_19             <= "000";
                soft_input_39                   <= (others => (others => '0'));
        elsif rising_edge(clk) then 
                soft_input_39                   <= soft_input_38;
                indi_4                          <= indi_3 and (corrections_temp_18 >= 0) and (corrections_temp_18 < 4); 
                hard_output_error_rest_21       <= hard_output_error_rest_20;                          -- pass the corrected data
                last_bit_1                      <= last_bit;                                           -- flip it anyway, store it here
                error_position_temp_19          <= error_position_temp_18;                             -- passing the error position
                corrections_temp_19             <= corrections_temp_18;                                -- passing the correction number
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 23)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then
                hard_output_error_rest_22                 <= (others => '0'); 
                error_position_temp_20(0)                 <= -1;
                error_position_temp_20(1)                 <= -1;
                error_position_temp_20(2)                 <= -1;
                corrections_temp_20                       <= "000";   
                soft_input_40                             <= (others => (others => '0'));  
        elsif rising_edge(clk) then 
                soft_input_40                             <= soft_input_39;
                if indi_4 then                                  -- The last bit is wrong, correct it
                        hard_output_error_rest_22         <= hard_output_error_rest_21;
                        hard_output_error_rest_22(255)    <= last_bit_1;
                        error_position_temp_20            <= error_position_temp_19;
                        error_position_temp_20(2)         <= 256;
                        corrections_temp_20               <= corrections_temp_19 + "001";
                else                                            -- The last bit is okay, pass the data
                        hard_output_error_rest_22         <= hard_output_error_rest_21;
                        error_position_temp_20            <= error_position_temp_19;
                        corrections_temp_20               <= corrections_temp_19;
                end if;
        end if;
end process;
--------------------------------------------------------------------------------------------------------------
---- Define processes : (CLK 24)
--------------------------------------------------------------------------------------------------------------
process(clk, reset)
begin
	if (reset = '1') then   
                hard_output       <= (others => '0');
                corrections       <= (others => '0');       
                error_position(0) <= -1;
                error_position(1) <= -1;
                error_position(2) <= -1;
                soft_output       <= (others => (others => '0')); 
        elsif rising_edge(clk) then 
                hard_output       <= hard_output_error_rest_22;
                corrections       <= corrections_temp_20;
                error_position    <= error_position_temp_20;
                soft_output       <= soft_input_40;
        end if; 
end process;
end architecture;