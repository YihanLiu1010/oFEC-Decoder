-- Dual-Port Block RAM with Two Write Ports
-- Correct Modelization with a Shared Variable
-- Size of this RAM should be 8960 rows * 1 column, each 256 rows contains 1 input_data_array
library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.arr_pkg_1.all;
use work.arr_pkg_2.all;
use work.arr_pkg_3.all;
use work.arr_pkg_4.all;
use work.arr_pkg_5.all;
use work.arr_pkg_6.all;
entity ram is
    port (
        addra : in std_logic_vector(8 downto 0); -- It goes up to 280
        addrb : in std_logic_vector(8 downto 0);
        clka  : in std_logic;
        clkb  : in std_logic;
        dia   : in std_logic_vector(2047 downto 0); -- IN / OUT will be 1 square
        dib   : in std_logic_vector(2047 downto 0);
        ena   : in std_logic;
        enb   : in std_logic;
        wea   : in std_logic;
        web   : in std_logic;
        doa   : out std_logic_vector(2047 downto 0);
        dob   : out std_logic_vector(2047 downto 0)
    );
end ram;

architecture rtl of ram is
    type ramtype is array(0 to 295) of std_logic_vector(2047 downto 0); -- 256*8
    signal A_0 : std_logic_vector(2047 downto 0) := ("00000000000000010000001000000011000001000000010100000110000001110000100000001001000010100000101100001100000011010000111000001111000100000001000100010010000100110001010000010101000101100001011100011000000110010001101000011011000111000001110100011110000111110010000000100001001000100010001100100100001001010010011000100111001010000010100100101010001010110010110000101101001011100010111100110000001100010011001000110011001101000011010100110110001101110011100000111001001110100011101100111100001111010011111000111111010000000100000101000010010000110100010001000101010001100100011101001000010010010100101001001011010011000100110101001110010011110101000001010001010100100101001101010100010101010101011001010111010110000101100101011010010110110101110001011101010111100101111101100000011000010110001001100011011001000110010101100110011001110110100001101001011010100110101101101100011011010110111001101111011100000111000101110010011100110111010001110101011101100111011101111000011110010111101001111011011111000111110101111110011111111000000010000001100000101000001110000100100001011000011010000111100010001000100110001010100010111000110010001101100011101000111110010000100100011001001010010011100101001001010110010110100101111001100010011001100110101001101110011100100111011001111010011111101000001010000110100010101000111010010010100101101001101010011110101000101010011010101010101011101011001010110110101110101011111011000010110001101100101011001110110100101101011011011010110111101110001011100110111010101110111011110010111101101111101011111111000000110000011100001011000011110001001100010111000110110001111100100011001001110010101100101111001100110011011100111011001111110100001101000111010010110100111101010011010101110101101101011111011000110110011101101011011011110111001101110111011110110111111110000011100001111000101110001111100100111001011110011011100111111010001110100111101010111010111110110011101101111011101110111111110000111100011111001011110011111101001111010111110110111101111111100011111001111110101111101111111100111111011111111011111111");
    signal A_1 : std_logic_vector(2047 downto 0) := ("00000001000000100000001100000100000001010000011000000111000010000000100100001010000010110000110000001101000011100000111100010000000100010001001000010011000101000001010100010110000101110001100000011001000110100001101100011100000111010001111000011111001000000010000100100010001000110010010000100101001001100010011100101000001010010010101000101011001011000010110100101110001011110011000000110001001100100011001100110100001101010011011000110111001110000011100100111010001110110011110000111101001111100011111101000000010000010100001001000011010001000100010101000110010001110100100001001001010010100100101101001100010011010100111001001111010100000101000101010010010100110101010001010101010101100101011101011000010110010101101001011011010111000101110101011110010111110110000001100001011000100110001101100100011001010110011001100111011010000110100101101010011010110110110001101101011011100110111101110000011100010111001001110011011101000111010101110110011101110111100001111001011110100111101101111100011111010111111001111111100000001000000110000010100000111000010010000101100001101000011110001000100010011000101010001011100011001000110110001110100011111001000010010001100100101001001110010100100101011001011010010111100110001001100110011010100110111001110010011101100111101001111110100000101000011010001010100011101001001010010110100110101001111010100010101001101010101010101110101100101011011010111010101111101100001011000110110010101100111011010010110101101101101011011110111000101110011011101010111011101111001011110110111110101111111100000011000001110000101100001111000100110001011100011011000111110010001100100111001010110010111100110011001101110011101100111111010000110100011101001011010011110101001101010111010110110101111101100011011001110110101101101111011100110111011101111011011111111000001110000111100010111000111110010011100101111001101110011111101000111010011110101011101011111011001110110111101110111011111111000011110001111100101111001111110100111101011111011011110111111110001111100111111010111110111111110011111101111111101111111100000000");
    signal A_2 : std_logic_vector(2047 downto 0) := ("00000010000000110000010000000101000001100000011100001000000010010000101000001011000011000000110100001110000011110001000000010001000100100001001100010100000101010001011000010111000110000001100100011010000110110001110000011101000111100001111100100000001000010010001000100011001001000010010100100110001001110010100000101001001010100010101100101100001011010010111000101111001100000011000100110010001100110011010000110101001101100011011100111000001110010011101000111011001111000011110100111110001111110100000001000001010000100100001101000100010001010100011001000111010010000100100101001010010010110100110001001101010011100100111101010000010100010101001001010011010101000101010101010110010101110101100001011001010110100101101101011100010111010101111001011111011000000110000101100010011000110110010001100101011001100110011101101000011010010110101001101011011011000110110101101110011011110111000001110001011100100111001101110100011101010111011001110111011110000111100101111010011110110111110001111101011111100111111110000000100000011000001010000011100001001000010110000110100001111000100010001001100010101000101110001100100011011000111010001111100100001001000110010010100100111001010010010101100101101001011110011000100110011001101010011011100111001001110110011110100111111010000010100001101000101010001110100100101001011010011010100111101010001010100110101010101010111010110010101101101011101010111110110000101100011011001010110011101101001011010110110110101101111011100010111001101110101011101110111100101111011011111010111111110000001100000111000010110000111100010011000101110001101100011111001000110010011100101011001011110011001100110111001110110011111101000011010001110100101101001111010100110101011101011011010111110110001101100111011010110110111101110011011101110111101101111111100000111000011110001011100011111001001110010111100110111001111110100011101001111010101110101111101100111011011110111011101111111100001111000111110010111100111111010011110101111101101111011111111000111110011111101011111011111111001111110111111110111111110000000000000001");
    signal A_3 : std_logic_vector(2047 downto 0) := ("00000011000001000000010100000110000001110000100000001001000010100000101100001100000011010000111000001111000100000001000100010010000100110001010000010101000101100001011100011000000110010001101000011011000111000001110100011110000111110010000000100001001000100010001100100100001001010010011000100111001010000010100100101010001010110010110000101101001011100010111100110000001100010011001000110011001101000011010100110110001101110011100000111001001110100011101100111100001111010011111000111111010000000100000101000010010000110100010001000101010001100100011101001000010010010100101001001011010011000100110101001110010011110101000001010001010100100101001101010100010101010101011001010111010110000101100101011010010110110101110001011101010111100101111101100000011000010110001001100011011001000110010101100110011001110110100001101001011010100110101101101100011011010110111001101111011100000111000101110010011100110111010001110101011101100111011101111000011110010111101001111011011111000111110101111110011111111000000010000001100000101000001110000100100001011000011010000111100010001000100110001010100010111000110010001101100011101000111110010000100100011001001010010011100101001001010110010110100101111001100010011001100110101001101110011100100111011001111010011111101000001010000110100010101000111010010010100101101001101010011110101000101010011010101010101011101011001010110110101110101011111011000010110001101100101011001110110100101101011011011010110111101110001011100110111010101110111011110010111101101111101011111111000000110000011100001011000011110001001100010111000110110001111100100011001001110010101100101111001100110011011100111011001111110100001101000111010010110100111101010011010101110101101101011111011000110110011101101011011011110111001101110111011110110111111110000011100001111000101110001111100100111001011110011011100111111010001110100111101010111010111110110011101101111011101110111111110000111100011111001011110011111101001111010111110110111101111111100011111001111110101111101111111100111111011111111011111111000000000000000100000010");
    signal A_4 : std_logic_vector(2047 downto 0) := ("00000100000001010000011000000111000010000000100100001010000010110000110000001101000011100000111100010000000100010001001000010011000101000001010100010110000101110001100000011001000110100001101100011100000111010001111000011111001000000010000100100010001000110010010000100101001001100010011100101000001010010010101000101011001011000010110100101110001011110011000000110001001100100011001100110100001101010011011000110111001110000011100100111010001110110011110000111101001111100011111101000000010000010100001001000011010001000100010101000110010001110100100001001001010010100100101101001100010011010100111001001111010100000101000101010010010100110101010001010101010101100101011101011000010110010101101001011011010111000101110101011110010111110110000001100001011000100110001101100100011001010110011001100111011010000110100101101010011010110110110001101101011011100110111101110000011100010111001001110011011101000111010101110110011101110111100001111001011110100111101101111100011111010111111001111111100000001000000110000010100000111000010010000101100001101000011110001000100010011000101010001011100011001000110110001110100011111001000010010001100100101001001110010100100101011001011010010111100110001001100110011010100110111001110010011101100111101001111110100000101000011010001010100011101001001010010110100110101001111010100010101001101010101010101110101100101011011010111010101111101100001011000110110010101100111011010010110101101101101011011110111000101110011011101010111011101111001011110110111110101111111100000011000001110000101100001111000100110001011100011011000111110010001100100111001010110010111100110011001101110011101100111111010000110100011101001011010011110101001101010111010110110101111101100011011001110110101101101111011100110111011101111011011111111000001110000111100010111000111110010011100101111001101110011111101000111010011110101011101011111011001110110111101110111011111111000011110001111100101111001111110100111101011111011011110111111110001111100111111010111110111111110011111101111111101111111100000000000000010000001000000011");
    --signal A_5 : std_logic_vector(2047 downto 0) := ("00000101000001100000011100001000000010010000101000001011000011000000110100001110000011110001000000010001000100100001001100010100000101010001011000010111000110000001100100011010000110110001110000011101000111100001111100100000001000010010001000100011001001000010010100100110001001110010100000101001001010100010101100101100001011010010111000101111001100000011000100110010001100110011010000110101001101100011011100111000001110010011101000111011001111000011110100111110001111110100000001000001010000100100001101000100010001010100011001000111010010000100100101001010010010110100110001001101010011100100111101010000010100010101001001010011010101000101010101010110010101110101100001011001010110100101101101011100010111010101111001011111011000000110000101100010011000110110010001100101011001100110011101101000011010010110101001101011011011000110110101101110011011110111000001110001011100100111001101110100011101010111011001110111011110000111100101111010011110110111110001111101011111100111111110000000100000011000001010000011100001001000010110000110100001111000100010001001100010101000101110001100100011011000111010001111100100001001000110010010100100111001010010010101100101101001011110011000100110011001101010011011100111001001110110011110100111111010000010100001101000101010001110100100101001011010011010100111101010001010100110101010101010111010110010101101101011101010111110110000101100011011001010110011101101001011010110110110101101111011100010111001101110101011101110111100101111011011111010111111110000001100000111000010110000111100010011000101110001101100011111001000110010011100101011001011110011001100110111001110110011111101000011010001110100101101001111010100110101011101011011010111110110001101100111011010110110111101110011011101110111101101111111100000111000011110001011100011111001001110010111100110111001111110100011101001111010101110101111101100111011011110111011101111111100001111000111110010111100111111010011110101111101101111011111111000111110011111101011111011111111001111110111111110111111110000000000000001000000100000001100000100");

    shared variable RAM : ramtype := (A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4,
    A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4,
    A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4,
    A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4,
    A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4,
    A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4,
    A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0, A_1, A_2, A_3, A_4, A_0);
begin

    process (CLKA)
    begin
        if CLKA'event and CLKA = '1' then
            if ENA = '1' then
                DOA <= RAM(to_integer(unsigned(ADDRA)));
                if WEA = '1' then
                    RAM(to_integer(unsigned(ADDRA))) := DIA;
                end if;
            end if;
        end if;
    end process;

    process (CLKB)
    begin
        if CLKB'event and CLKB = '1' then
            if ENB = '1' then
                DOB <= RAM(to_integer(unsigned(ADDRB)));
                if WEB = '1' then
                    RAM(to_integer(unsigned(ADDRB))) := DIB;
                end if;
            end if;
        end if;
    end process;
end architecture;
