library ieee;
use STD.textio.all;
use ieee.std_logic_textio.all;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use work.arr_pkg_1.all;
use work.arr_pkg_2.all;
use work.arr_pkg_3.all;
use work.arr_pkg_4.all;
use work.arr_pkg_5.all;
use work.arr_pkg_6.all;
-- Seperation for writing data back should be done in Extrinsic calculation!!! Otherwise there might not be enough time
entity ram_top is
    port (
        clk   : in std_logic;
        reset : in std_logic;
        -- Write data back, put all 16 codewords together(16*256)
        -- dat_i : in input_data_array(4095 downto 0);
        data_in_1 : in std_logic_vector(2047 downto 0);
        data_in_2 : in std_logic_vector(2047 downto 0);
        rdreq     : in std_logic;
        wrreq     : in std_logic;
        -- Read data out, I only need half, the other half comes from the channel
        --dat_o : out input_data_array(2047 downto 0)
        data_out_1 : out std_logic_vector(2047 downto 0);
        data_out_2 : out std_logic_vector(2047 downto 0)
    );
end ram_top;
architecture rtl of ram_top is
    -----------------------------------------------------------------------------------------------------------
    -- pre-calcaulated array
    type table_1 is array (0 to 296) of std_logic_vector(8 downto 0); -- Read address table
    type table_2 is array (0 to 591) of std_logic_vector(8 downto 0); -- Write address table
    constant addr_table_1 : table_1 := (
        "011101000","011110001","011111010","100000011","100001100","100010101","100011110","100100111",
        "011110000","011111001","100000010","100001011","100010100","100011101","100100110","000000111",
        "011111000","100000001","100001010","100010011","100011100","100100101","000000110","000001111",
        "100000000","100001001","100010010","100011011","100100100","000000101","000001110","000010111",
        "100001000","100010001","100011010","100100011","000000100","000001101","000010110","000011111",
        "100010000","100011001","100100010","000000011","000001100","000010101","000011110","000100111",
        "100011000","100100001","000000010","000001011","000010100","000011101","000100110","000101111",
        "100100000","000000001","000001010","000010011","000011100","000100101","000101110","000110111",
        "000000000","000001001","000010010","000011011","000100100","000101101","000110110","000111111",
        "000001000","000010001","000011010","000100011","000101100","000110101","000111110","001000111",
        "000010000","000011001","000100010","000101011","000110100","000111101","001000110","001001111",
        "000011000","000100001","000101010","000110011","000111100","001000101","001001110","001010111",
        "000100000","000101001","000110010","000111011","001000100","001001101","001010110","001011111",
        "000101000","000110001","000111010","001000011","001001100","001010101","001011110","001100111",
        "000110000","000111001","001000010","001001011","001010100","001011101","001100110","001101111",
        "000111000","001000001","001001010","001010011","001011100","001100101","001101110","001110111",
        "001000000","001001001","001010010","001011011","001100100","001101101","001110110","001111111",
        "001001000","001010001","001011010","001100011","001101100","001110101","001111110","010000111",
        "001010000","001011001","001100010","001101011","001110100","001111101","010000110","010001111",
        "001011000","001100001","001101010","001110011","001111100","010000101","010001110","010010111",
        "001100000","001101001","001110010","001111011","010000100","010001101","010010110","010011111",
        "001101000","001110001","001111010","010000011","010001100","010010101","010011110","010100111",
        "001110000","001111001","010000010","010001011","010010100","010011101","010100110","010101111",
        "001111000","010000001","010001010","010010011","010011100","010100101","010101110","010110111",
        "010000000","010001001","010010010","010011011","010100100","010101101","010110110","010111111",
        "010001000","010010001","010011010","010100011","010101100","010110101","010111110","011000111",
        "010010000","010011001","010100010","010101011","010110100","010111101","011000110","011001111",
        "010011000","010100001","010101010","010110011","010111100","011000101","011001110","011010111",
        "010100000","010101001","010110010","010111011","011000100","011001101","011010110","011011111",
        "010101000","010110001","010111010","011000011","011001100","011010101","011011110","011100111",
        "010110000","010111001","011000010","011001011","011010100","011011101","011100110","011101111",
        "010111000","011000001","011001010","011010011","011011100","011100101","011101110","011110111",
        "011000000","011001001","011010010","011011011","011100100","011101101","011110110","011111111",
        "011001000","011010001","011011010","011100011","011101100","011110101","011111110","100000111",
        "011010000","011011001","011100010","011101011","011110100","011111101","100000110","100001111",
        "011011000","011100001","011101010","011110011","011111100","100000101","100001110","100010111",
        "011100000","011101001","011110010","011111011","100000100","100001101","100010110","100011111", "111111111"
    );
    constant addr_table_3 : table_2 := (
        "001101000", "001110001", "001111010", "010000011", "010001100", "010010101", "010011110", "010100111", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
        "001110000", "001111001", "010000010", "010001011", "010010100", "010011101", "010100110", "010101111", "000000001", "000000001", "000000001", "000000001", "000000001", "000000001", "000000001", "000000001",
        "001111000", "010000001", "010001010", "010010011", "010011100", "010100101", "010101110", "010110111", "000000010", "000000010", "000000010", "000000010", "000000010", "000000010", "000000010", "000000010",
        "010000000", "010001001", "010010010", "010011011", "010100100", "010101101", "010110110", "010111111", "000000011", "000000011", "000000011", "000000011", "000000011", "000000011", "000000011", "000000011",
        "010001000", "010010001", "010011010", "010100011", "010101100", "010110101", "010111110", "011000111", "000000100", "000000100", "000000100", "000000100", "000000100", "000000100", "000000100", "000000100",
        "010010000", "010011001", "010100010", "010101011", "010110100", "010111101", "011000110", "011001111", "000000101", "000000101", "000000101", "000000101", "000000101", "000000101", "000000101", "000000101",
        "010011000", "010100001", "010101010", "010110011", "010111100", "011000101", "011001110", "011010111", "000000110", "000000110", "000000110", "000000110", "000000110", "000000110", "000000110", "000000110",
        "010100000", "010101001", "010110010", "010111011", "011000100", "011001101", "011010110", "011011111", "000000111", "000000111", "000000111", "000000111", "000000111", "000000111", "000000111", "000000111",
        "010101000", "010110001", "010111010", "011000011", "011001100", "011010101", "011011110", "011100111", "000001000", "000001000", "000001000", "000001000", "000001000", "000001000", "000001000", "000001000",
        "010110000", "010111001", "011000010", "011001011", "011010100", "011011101", "011100110", "011101111", "000001001", "000001001", "000001001", "000001001", "000001001", "000001001", "000001001", "000001001",
        "010111000", "011000001", "011001010", "011010011", "011011100", "011100101", "011101110", "011110111", "000001010", "000001010", "000001010", "000001010", "000001010", "000001010", "000001010", "000001010",
        "011000000", "011001001", "011010010", "011011011", "011100100", "011101101", "011110110", "011111111", "000001011", "000001011", "000001011", "000001011", "000001011", "000001011", "000001011", "000001011",
        "011001000", "011010001", "011011010", "011100011", "011101100", "011110101", "011111110", "100000111", "000001100", "000001100", "000001100", "000001100", "000001100", "000001100", "000001100", "000001100",
        "011010000", "011011001", "011100010", "011101011", "011110100", "011111101", "100000110", "100001111", "000001101", "000001101", "000001101", "000001101", "000001101", "000001101", "000001101", "000001101",
        "011011000", "011100001", "011101010", "011110011", "011111100", "100000101", "100001110", "100010111", "000001110", "000001110", "000001110", "000001110", "000001110", "000001110", "000001110", "000001110",
        "011100000", "011101001", "011110010", "011111011", "100000100", "100001101", "100010110", "000000111", "000001111", "000001111", "000001111", "000001111", "000001111", "000001111", "000001111", "000001111",
        "011101000", "011110001", "011111010", "100000011", "100001100", "100010101", "000000110", "000001111", "000010000", "000010000", "000010000", "000010000", "000010000", "000010000", "000010000", "000010000",
        "011110000", "011111001", "100000010", "100001011", "100010100", "000000101", "000001110", "000010111", "000010001", "000010001", "000010001", "000010001", "000010001", "000010001", "000010001", "000010001",
        "011111000", "100000001", "100001010", "100010011", "000000100", "000001101", "000010110", "000011111", "000010010", "000010010", "000010010", "000010010", "000010010", "000010010", "000010010", "000010010",
        "100000000", "100001001", "100010010", "000000011", "000001100", "000010101", "000011110", "000100111", "000010011", "000010011", "000010011", "000010011", "000010011", "000010011", "000010011", "000010011",
        "100001000", "100010001", "000000010", "000001011", "000010100", "000011101", "000100110", "000101111", "000010100", "000010100", "000010100", "000010100", "000010100", "000010100", "000010100", "000010100",
        "100010000", "000000001", "000001010", "000010011", "000011100", "000100101", "000101110", "000110111", "000010101", "000010101", "000010101", "000010101", "000010101", "000010101", "000010101", "000010101",
        "000000000", "000001001", "000010010", "000011011", "000100100", "000101101", "000110110", "000111111", "000010110", "000010110", "000010110", "000010110", "000010110", "000010110", "000010110", "000010110",
        "000001000", "000010001", "000011010", "000100011", "000101100", "000110101", "000111110", "001000111", "000010111", "000010111", "000010111", "000010111", "000010111", "000010111", "000010111", "000010111",
        "000010000", "000011001", "000100010", "000101011", "000110100", "000111101", "001000110", "001001111", "000011000", "000011000", "000011000", "000011000", "000011000", "000011000", "000011000", "000011000",
        "000011000", "000100001", "000101010", "000110011", "000111100", "001000101", "001001110", "001010111", "000011001", "000011001", "000011001", "000011001", "000011001", "000011001", "000011001", "000011001",
        "000100000", "000101001", "000110010", "000111011", "001000100", "001001101", "001010110", "001011111", "000011010", "000011010", "000011010", "000011010", "000011010", "000011010", "000011010", "000011010",
        "000101000", "000110001", "000111010", "001000011", "001001100", "001010101", "001011110", "001100111", "000011011", "000011011", "000011011", "000011011", "000011011", "000011011", "000011011", "000011011",
        "000110000", "000111001", "001000010", "001001011", "001010100", "001011101", "001100110", "001101111", "000011100", "000011100", "000011100", "000011100", "000011100", "000011100", "000011100", "000011100",
        "000111000", "001000001", "001001010", "001010011", "001011100", "001100101", "001101110", "001110111", "000011101", "000011101", "000011101", "000011101", "000011101", "000011101", "000011101", "000011101",
        "001000000", "001001001", "001010010", "001011011", "001100100", "001101101", "001110110", "001111111", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110",
        "001001000", "001010001", "001011010", "001100011", "001101100", "001110101", "001111110", "010000111", "000011111", "000011111", "000011111", "000011111", "000011111", "000011111", "000011111", "000011111",
        "001010000", "001011001", "001100010", "001101011", "001110100", "001111101", "010000110", "010001111", "000100000", "000100000", "000100000", "000100000", "000100000", "000100000", "000100000", "000100000",
        "001011000", "001100001", "001101010", "001110011", "001111100", "010000101", "010001110", "010010111", "000100001", "000100001", "000100001", "000100001", "000100001", "000100001", "000100001", "000100001",
        "001100000", "001101001", "001110010", "001111011", "010000100", "010001101", "010010110", "010011111", "000100010", "000100010", "000100010", "000100010", "000100010", "000100010", "000100010", "000100010",
        "001011000", "001100001", "001101010", "001110011", "001111100", "010000101", "010001110", "010010111", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011",
        "001100000", "001101001", "001110010", "001111011", "010000100", "010001101", "010010110", "010011111", "000100100", "000100100", "000100100", "000100100", "000100100", "000100100", "000100100", "000100100"
    );
    signal rdreq_a_1, rdreq_a_2, wrreq_a_1, wrreq_a_2               : std_logic;
    signal addr_write                                               : std_logic_vector(8 downto 0);
    signal addr_a_read_1, addr_a_read_2, addr_a_1, addr_a_2         : std_logic_vector(8 downto 0);
    signal q_a_1, q_a_2, data_a_1, data_a_2, data_a_1_r, data_a_2_r : std_logic_vector(2047 downto 0);
    signal i                                                        : std_logic_vector(9 downto 0) := (others => '0');
    signal j                                                        : integer range 0 to 296;
    signal output_index                                             : integer := 0;

begin

    ram_a : entity work.ram port map(addr_a_1, addr_a_2, clk, clk, data_a_1, data_a_2, rdreq_a_1, rdreq_a_2, wrreq_a_1, wrreq_a_2, q_a_1, q_a_2);

    data_out_1 <= q_a_1; -- output
    data_out_2 <= q_a_2;
    data_a_1   <= data_in_1;--input
    data_a_2   <= data_in_2;

    trans : process (clk)
    begin
        if (reset = '1') then
            addr_a_read_1 <= (others => '0');
            addr_a_read_2 <= (others => '0');
            i             <= (others => '0');
            data_a_1      <= (others => '0');
            data_a_2      <= (others => '0');
        else
            if (rising_edge(clk)) then
                if (rdreq = '1') then -- Get the reading done!
                    if i(0) = '0' then    -- even number
                        addr_a_1 <= addr_table_1(0 + j);
                        j        <= j + 1;
                    else
                        addr_a_1 <= addr_a_1;
                        j        <= j;
                    end if;
                    rdreq_a_1 <= '1'; -- Read request
                    if (i = "1001001111") then
                        i <= "0000000000";
                        j <= 0;
                    else
                        i <= i + '1';
                    end if;
                else
                    rdreq_a_1 <= '0';
                end if;
                if (wrreq = '1') then -- writing back is also half speed
                    wrreq_a_1 <= '1';     -- write request
                    wrreq_a_2 <= '1';
                    addr_a_1  <= addr_write;
                    addr_a_2  <= addr_write + 1;
                    data_a_1  <= data_a_1_r;
                    data_a_2  <= data_a_2_r;
                else
                    wrreq_a_1 <= '0';
                    wrreq_a_2 <= '0';
                end if;
            end if;
        end if;
    end process;
end architecture;
